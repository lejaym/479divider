magic
tech scmos
timestamp 1428359926
<< pwell >>
rect 903 1221 910 1234
<< metal1 >>
rect -34 1749 4 1822
rect 910 1807 976 1823
rect -34 1733 30 1749
rect -34 1560 4 1733
rect 938 1675 976 1807
rect 909 1659 976 1675
rect 915 1635 920 1643
rect 910 1617 920 1623
rect -34 1544 30 1560
rect -34 1359 4 1544
rect 910 1446 919 1454
rect 938 1433 976 1659
rect 910 1417 976 1433
rect -34 1339 30 1359
rect -34 1124 4 1339
rect 938 1320 976 1417
rect 910 1316 976 1320
rect 938 1229 976 1316
rect 910 1221 976 1229
rect -34 1116 30 1124
rect -34 893 4 1116
rect 938 1021 976 1221
rect 938 998 1865 1021
rect 910 997 1865 998
rect 909 993 1865 997
rect 1785 986 1865 993
rect -34 878 30 893
rect -34 670 4 878
rect 1795 745 1807 753
rect 1790 727 1807 733
rect -34 654 30 670
rect -34 524 4 654
rect 1828 555 1865 986
rect 1790 547 1865 555
rect -34 513 30 524
rect -34 385 4 513
rect -34 369 30 385
rect -34 237 4 369
rect 1828 311 1865 547
rect 1790 295 1865 311
rect 1790 267 1798 277
rect -34 220 30 237
rect -34 36 4 220
rect 1790 123 1798 131
rect 1828 110 1865 295
rect 1790 94 1865 110
rect -34 20 31 36
rect 1828 19 1865 94
<< metal2 >>
rect 43 1823 49 1864
rect 153 1823 159 1864
rect 263 1823 269 1864
rect 373 1823 379 1864
rect 483 1823 489 1864
rect 593 1823 599 1864
rect 703 1823 709 1864
rect 813 1823 819 1864
rect 1005 994 1011 1073
rect 1115 994 1121 1073
rect 1225 994 1231 1073
rect 1335 994 1341 1073
rect 1445 994 1451 1073
rect 1555 994 1561 1073
rect 1665 994 1671 1073
rect 1774 994 1780 1073
rect 1790 493 1815 501
rect 1790 466 1814 469
rect 1794 462 1814 466
rect 81 -21 94 20
rect 191 -21 204 20
rect 301 -21 314 20
rect 411 -21 424 20
rect 521 -21 534 20
rect 631 -21 644 20
rect 741 -21 754 20
rect 851 -21 864 20
rect 961 -21 974 20
rect 1071 -21 1084 20
rect 1181 -21 1194 20
rect 1291 -21 1304 20
rect 1401 -21 1414 20
rect 1511 -21 1524 20
rect 1621 -21 1634 20
rect 1731 -21 1744 20
<< polycontact >>
rect 910 1635 915 1643
rect 1790 745 1795 753
<< m2contact >>
rect 920 1635 925 1643
rect 920 1617 925 1623
rect 919 1446 925 1454
rect 1807 745 1812 753
rect 1807 727 1812 733
rect 1790 462 1794 466
rect 1798 267 1806 277
rect 1798 123 1804 131
use datapathL  datapathL_0 ../cells
array 0 7 110 0 0 1803
timestamp 1428357410
transform 1 0 30 0 1 562
box 0 -542 110 1261
use datapathS  datapathS_0 ../cells
array 0 7 110 0 0 974
timestamp 1428358217
transform 1 0 910 0 1 562
box 0 -542 110 432
<< labels >>
rlabel metal2 1790 495 1815 499 0 INBIT
rlabel metal1 -34 20 4 1822 0 Vdd
rlabel metal1 1828 19 1865 1021 0 GND
<< end >>
