magic
tech scmos
timestamp 1428347008
<< pwell >>
rect -49 113 -26 142
rect -49 73 41 113
rect -49 -42 41 -2
rect -49 -71 -26 -42
<< nwell >>
rect -23 117 41 147
rect -49 2 41 69
rect -22 -76 41 -46
<< polysilicon >>
rect -36 141 -23 143
rect -36 140 -34 141
rect -25 140 -23 141
rect -12 138 -10 149
rect -2 138 0 150
rect 8 138 10 140
rect 18 138 20 140
rect -12 110 -10 120
rect -2 110 0 120
rect 8 117 10 120
rect 18 118 20 120
rect 8 113 9 117
rect 18 114 29 118
rect 8 110 10 113
rect 18 110 20 114
rect -36 98 -34 100
rect -30 88 -19 90
rect -40 86 -38 88
rect -30 86 -28 88
rect -40 66 -38 76
rect -30 66 -28 76
rect -21 69 -19 88
rect -12 86 -10 100
rect -2 86 0 100
rect 8 98 10 100
rect 18 98 20 100
rect 8 86 10 88
rect 18 86 20 88
rect -12 66 -10 76
rect -2 74 0 76
rect 8 74 10 76
rect -2 72 10 74
rect -2 66 0 72
rect 8 66 10 72
rect 18 66 20 76
rect -40 32 -38 46
rect -30 44 -28 46
rect -12 32 -10 46
rect -40 28 -39 32
rect -11 28 -10 32
rect -40 25 -38 28
rect -22 25 -20 27
rect -12 25 -10 28
rect -2 32 0 46
rect 8 44 10 46
rect 18 40 20 46
rect 18 38 28 40
rect 26 32 28 38
rect -2 28 -1 32
rect 27 28 28 32
rect -2 25 0 28
rect 8 25 10 27
rect 26 25 28 28
rect -40 -5 -38 5
rect -22 2 -20 5
rect -31 -2 -20 2
rect -22 -5 -20 -2
rect -12 -5 -10 5
rect -2 -5 0 5
rect 8 2 10 5
rect 8 -2 19 2
rect 8 -5 10 -2
rect 26 -5 28 5
rect -40 -17 -38 -15
rect -22 -17 -20 -15
rect -36 -29 -34 -27
rect -12 -29 -10 -15
rect -2 -29 0 -15
rect 8 -17 10 -15
rect 26 -17 28 -15
rect 8 -29 10 -27
rect -12 -49 -10 -39
rect -2 -49 0 -39
rect 8 -42 10 -39
rect 8 -46 9 -42
rect 8 -49 10 -46
rect -36 -70 -34 -69
rect -25 -70 -23 -69
rect -36 -72 -23 -70
rect -12 -79 -10 -67
rect -2 -79 0 -67
rect 8 -81 10 -67
<< ndiffusion >>
rect -38 100 -36 140
rect -34 100 -32 140
rect -14 100 -12 110
rect -10 100 -2 110
rect 0 100 8 110
rect 10 100 12 110
rect 16 100 18 110
rect 20 100 22 110
rect -42 76 -40 86
rect -38 76 -36 86
rect -32 76 -30 86
rect -28 76 -26 86
rect -14 76 -12 86
rect -10 76 -8 86
rect -4 76 -2 86
rect 0 76 2 86
rect 6 76 8 86
rect 10 76 18 86
rect 20 76 22 86
rect -42 -15 -40 -5
rect -38 -15 -36 -5
rect -24 -15 -22 -5
rect -20 -15 -18 -5
rect -14 -15 -12 -5
rect -10 -15 -8 -5
rect -4 -15 -2 -5
rect 0 -15 2 -5
rect 6 -15 8 -5
rect 10 -15 12 -5
rect 24 -15 26 -5
rect 28 -15 30 -5
rect -38 -69 -36 -29
rect -34 -69 -32 -29
rect -14 -39 -12 -29
rect -10 -39 -2 -29
rect 0 -39 8 -29
rect 10 -39 12 -29
<< pdiffusion >>
rect -14 120 -12 138
rect -10 120 -8 138
rect -4 120 -2 138
rect 0 120 2 138
rect 6 120 8 138
rect 10 120 12 138
rect 16 120 18 138
rect 20 120 22 138
rect -42 46 -40 66
rect -38 46 -36 66
rect -32 46 -30 66
rect -28 46 -26 66
rect -14 46 -12 66
rect -10 46 -2 66
rect 0 46 2 66
rect 6 46 8 66
rect 10 46 12 66
rect 16 46 18 66
rect 20 46 22 66
rect -42 5 -40 25
rect -38 5 -36 25
rect -24 5 -22 25
rect -20 5 -18 25
rect -14 5 -12 25
rect -10 5 -8 25
rect -4 5 -2 25
rect 0 5 2 25
rect 6 5 8 25
rect 10 5 12 25
rect 24 5 26 25
rect 28 5 30 25
rect -14 -67 -12 -49
rect -10 -67 -8 -49
rect -4 -67 -2 -49
rect 0 -67 2 -49
rect 6 -67 8 -49
rect 10 -67 12 -49
<< metal1 >>
rect -60 143 30 147
rect -60 43 -53 143
rect -49 127 -45 131
rect -49 116 -45 120
rect -49 104 -45 108
rect -8 138 -4 143
rect 12 138 16 143
rect 40 143 41 147
rect -25 135 -21 136
rect -28 120 -18 125
rect -28 117 -14 120
rect 2 117 6 120
rect 22 117 26 120
rect -28 116 6 117
rect -28 112 -18 116
rect -14 113 6 116
rect 13 113 26 117
rect -28 110 -14 112
rect 22 110 26 113
rect -28 100 -18 110
rect 29 113 33 114
rect -42 97 -38 100
rect 12 97 16 100
rect -49 96 52 97
rect -49 90 -45 96
rect -31 90 6 96
rect 29 90 52 96
rect -49 89 52 90
rect -36 86 -32 89
rect -18 86 -14 89
rect 2 86 6 89
rect -46 73 -42 76
rect -49 69 -42 73
rect -46 66 -42 69
rect -26 73 -22 76
rect -8 73 -4 76
rect 22 73 26 76
rect -15 69 -8 73
rect 16 69 26 73
rect -26 66 -22 69
rect -18 66 -14 69
rect 12 66 16 69
rect -36 43 -32 46
rect 2 43 6 46
rect 22 43 26 46
rect -60 42 41 43
rect -60 35 -37 42
rect -16 35 41 42
rect -60 -72 -53 35
rect -46 25 -42 35
rect -35 28 -34 32
rect -16 28 -15 32
rect -8 25 -4 35
rect 3 28 4 32
rect 22 28 23 32
rect 30 25 34 35
rect -32 5 -31 25
rect -35 2 -31 5
rect -49 -2 -46 2
rect -28 2 -24 5
rect 12 2 16 5
rect -28 -2 -18 2
rect -35 -5 -31 -2
rect -18 -5 -14 -2
rect 6 -2 16 2
rect 19 5 20 25
rect 19 2 23 5
rect 2 -5 6 -2
rect 19 -5 23 -2
rect -32 -15 -31 -5
rect 19 -15 20 -5
rect -46 -18 -42 -15
rect -28 -18 -24 -15
rect -8 -18 -4 -15
rect 12 -18 16 -15
rect 30 -18 34 -15
rect 46 -18 52 89
rect -49 -19 52 -18
rect -49 -25 6 -19
rect 31 -25 52 -19
rect -49 -26 52 -25
rect -42 -29 -38 -26
rect 12 -29 16 -26
rect -49 -37 -45 -33
rect -49 -50 -45 -46
rect -28 -39 -18 -29
rect -28 -42 -14 -39
rect -28 -46 -18 -42
rect -14 -46 6 -42
rect 13 -46 29 -42
rect -28 -49 -14 -46
rect 2 -49 6 -46
rect -25 -65 -21 -64
rect -8 -72 -4 -67
rect 12 -72 16 -67
rect -60 -76 20 -72
rect 39 -76 41 -72
<< metal2 >>
rect -21 131 41 132
rect -25 128 41 131
rect -45 124 -38 127
rect -45 123 16 124
rect -42 120 16 123
rect -45 112 -18 116
rect -45 100 -4 104
rect -8 73 -4 100
rect 12 73 16 120
rect -49 65 -22 69
rect -20 36 22 40
rect -20 32 -16 36
rect 18 32 22 36
rect -34 24 -30 28
rect 4 24 8 28
rect -34 20 8 24
rect -42 -2 -18 2
rect 2 -29 6 -2
rect -45 -33 6 -29
rect 29 -42 33 109
rect -45 -46 -18 -42
rect 37 -50 41 128
rect -25 -54 41 -50
rect -25 -60 -21 -54
<< ntransistor >>
rect -36 100 -34 140
rect -12 100 -10 110
rect -2 100 0 110
rect 8 100 10 110
rect 18 100 20 110
rect -40 76 -38 86
rect -30 76 -28 86
rect -12 76 -10 86
rect -2 76 0 86
rect 8 76 10 86
rect 18 76 20 86
rect -40 -15 -38 -5
rect -22 -15 -20 -5
rect -12 -15 -10 -5
rect -2 -15 0 -5
rect 8 -15 10 -5
rect 26 -15 28 -5
rect -36 -69 -34 -29
rect -12 -39 -10 -29
rect -2 -39 0 -29
rect 8 -39 10 -29
<< ptransistor >>
rect -12 120 -10 138
rect -2 120 0 138
rect 8 120 10 138
rect 18 120 20 138
rect -40 46 -38 66
rect -30 46 -28 66
rect -12 46 -10 66
rect -2 46 0 66
rect 8 46 10 66
rect 18 46 20 66
rect -40 5 -38 25
rect -22 5 -20 25
rect -12 5 -10 25
rect -2 5 0 25
rect 8 5 10 25
rect 26 5 28 25
rect -12 -67 -10 -49
rect -2 -67 0 -49
rect 8 -67 10 -49
<< polycontact >>
rect -25 136 -21 140
rect 9 113 13 117
rect 29 114 33 118
rect -19 69 -15 73
rect -39 28 -35 32
rect -15 28 -11 32
rect -1 28 3 32
rect 23 28 27 32
rect -35 -2 -31 2
rect 19 -2 23 2
rect 9 -46 13 -42
rect -25 -69 -21 -65
<< ndcontact >>
rect -42 100 -38 140
rect -32 100 -28 140
rect -18 100 -14 110
rect 12 100 16 110
rect 22 100 26 110
rect -46 76 -42 86
rect -36 76 -32 86
rect -26 76 -22 86
rect -18 76 -14 86
rect -8 76 -4 86
rect 2 76 6 86
rect 22 76 26 86
rect -46 -15 -42 -5
rect -36 -15 -32 -5
rect -28 -15 -24 -5
rect -18 -15 -14 -5
rect -8 -15 -4 -5
rect 2 -15 6 -5
rect 12 -15 16 -5
rect 20 -15 24 -5
rect 30 -15 34 -5
rect -42 -69 -38 -29
rect -32 -69 -28 -29
rect -18 -39 -14 -29
rect 12 -39 16 -29
<< pdcontact >>
rect -18 120 -14 138
rect -8 120 -4 138
rect 2 120 6 138
rect 12 120 16 138
rect 22 120 26 138
rect -46 46 -42 66
rect -36 46 -32 66
rect -26 46 -22 66
rect -18 46 -14 66
rect 2 46 6 66
rect 12 46 16 66
rect 22 46 26 66
rect -46 5 -42 25
rect -36 5 -32 25
rect -28 5 -24 25
rect -18 5 -14 25
rect -8 5 -4 25
rect 2 5 6 25
rect 12 5 16 25
rect 20 5 24 25
rect 30 5 34 25
rect -18 -67 -14 -49
rect -8 -67 -4 -49
rect 2 -67 6 -49
rect 12 -67 16 -49
<< m2contact >>
rect -49 123 -45 127
rect -49 112 -45 116
rect -49 100 -45 104
rect -25 131 -21 135
rect -18 112 -14 116
rect 29 109 33 113
rect -26 69 -22 73
rect -8 69 -4 73
rect 12 69 16 73
rect -34 28 -30 32
rect -20 28 -16 32
rect 4 28 8 32
rect 18 28 22 32
rect -46 -2 -42 2
rect -18 -2 -14 2
rect 2 -2 6 2
rect -49 -33 -45 -29
rect -49 -46 -45 -42
rect -18 -46 -14 -42
rect 29 -46 33 -42
rect -25 -64 -21 -60
<< psubstratepcontact >>
rect -45 90 -31 96
rect 6 90 29 96
rect 6 -25 31 -19
<< nsubstratencontact >>
rect 30 140 40 147
rect -37 35 -16 42
rect 20 -76 39 -72
<< labels >>
rlabel metal1 -46 66 -42 76 1 sel1
rlabel metal2 -49 65 -22 69 1 sel0
rlabel metal1 -49 -2 -46 2 3 add
rlabel metal1 13 -46 29 -42 1 sign
rlabel polysilicon -2 -79 0 -69 1 SB0
rlabel polysilicon -12 -79 -10 -69 1 SB1
rlabel metal1 -60 -76 -53 147 3 Vdd
rlabel metal1 46 -26 52 97 7 Gnd
rlabel metal1 -18 113 6 117 1 nextSB0
rlabel metal1 -49 104 -45 108 1 load
rlabel metal1 -49 127 -45 131 1 shift
rlabel metal1 -49 -37 -45 -33 1 inbit
rlabel metal1 -18 -46 6 -42 1 nextSB1
rlabel metal2 -25 -54 41 -50 1 start
<< end >>
