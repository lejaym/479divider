magic
tech scmos
timestamp 1428889669
<< pwell >>
rect 0 191 110 278
rect 0 0 110 45
<< nwell >>
rect 0 282 110 349
rect 0 49 110 187
<< polysilicon >>
rect 64 342 66 344
rect 74 342 76 344
rect 44 305 46 308
rect 64 305 66 322
rect 74 319 76 322
rect 74 305 76 315
rect 44 275 46 285
rect 64 275 66 285
rect 74 275 76 285
rect 44 262 46 265
rect 64 255 66 265
rect 64 248 66 251
rect 74 248 76 265
rect 64 236 66 238
rect 74 236 76 238
rect 36 225 56 227
rect 36 224 40 225
rect 54 222 56 225
rect 64 222 66 224
rect 74 222 76 224
rect 54 211 56 212
rect 64 211 66 212
rect 54 209 66 211
rect 42 205 46 207
rect 44 204 46 205
rect 44 184 46 194
rect 44 162 46 164
rect 54 152 56 209
rect 64 204 66 206
rect 74 204 76 212
rect 74 200 77 204
rect 64 191 66 194
rect 64 184 66 187
rect 64 161 66 164
rect 64 152 66 154
rect 74 152 76 200
rect 54 132 56 133
rect 64 132 66 133
rect 44 130 66 132
rect 44 79 46 130
rect 55 110 56 113
rect 54 107 56 110
rect 64 110 65 113
rect 64 107 66 110
rect 43 75 46 79
rect 24 72 26 74
rect 34 72 36 74
rect 44 72 46 75
rect 54 72 56 87
rect 64 72 66 87
rect 74 72 76 133
rect 84 107 86 109
rect 84 57 86 87
rect 84 53 87 57
rect 24 49 26 52
rect 24 42 26 45
rect 34 42 36 52
rect 44 42 46 52
rect 54 42 56 52
rect 64 42 66 52
rect 74 49 76 52
rect 74 42 76 45
rect 24 30 26 32
rect 34 29 36 32
rect 44 30 46 32
rect 34 25 35 29
rect 54 17 56 32
rect 64 17 66 32
rect 74 30 76 32
rect 84 17 86 53
rect 54 5 56 7
rect 64 5 66 7
rect 84 5 86 7
<< ndiffusion >>
rect 42 265 44 275
rect 46 265 48 275
rect 62 265 64 275
rect 66 265 68 275
rect 72 265 74 275
rect 76 265 78 275
rect 62 238 64 248
rect 66 238 68 248
rect 72 238 74 248
rect 76 238 78 248
rect 52 212 54 222
rect 56 212 58 222
rect 62 212 64 222
rect 66 212 68 222
rect 72 212 74 222
rect 76 212 78 222
rect 42 194 44 204
rect 46 194 48 204
rect 62 194 64 204
rect 66 194 68 204
rect 22 32 24 42
rect 26 32 28 42
rect 32 32 34 42
rect 36 32 38 42
rect 42 32 44 42
rect 46 32 48 42
rect 52 32 54 42
rect 56 32 58 42
rect 62 32 64 42
rect 66 32 68 42
rect 72 32 74 42
rect 76 32 78 42
rect 52 7 54 17
rect 56 7 58 17
rect 62 7 64 17
rect 66 7 68 17
rect 82 7 84 17
rect 86 7 88 17
<< pdiffusion >>
rect 62 322 64 342
rect 66 322 68 342
rect 72 322 74 342
rect 76 322 78 342
rect 42 285 44 305
rect 46 285 48 305
rect 62 285 64 305
rect 66 285 68 305
rect 72 285 74 305
rect 76 285 78 305
rect 42 164 44 184
rect 46 164 48 184
rect 62 164 64 184
rect 66 164 68 184
rect 52 133 54 152
rect 56 133 58 152
rect 62 133 64 152
rect 66 133 68 152
rect 72 133 74 152
rect 76 133 78 152
rect 52 87 54 107
rect 56 87 58 107
rect 62 87 64 107
rect 66 87 68 107
rect 82 87 84 107
rect 86 87 88 107
rect 22 52 24 72
rect 26 52 28 72
rect 32 52 34 72
rect 36 52 38 72
rect 42 52 44 72
rect 46 52 48 72
rect 52 52 54 72
rect 56 52 58 72
rect 62 52 64 72
rect 66 52 68 72
rect 72 52 74 72
rect 76 52 78 72
<< metal1 >>
rect 0 345 110 349
rect 33 344 47 345
rect 33 340 43 344
rect 33 336 36 340
rect 40 336 43 340
rect 68 342 72 345
rect 0 322 53 326
rect 57 322 58 342
rect 82 322 83 342
rect 90 322 110 326
rect 90 319 94 322
rect 29 315 70 319
rect 77 315 94 319
rect 29 282 33 315
rect 66 312 70 315
rect 47 308 62 312
rect 66 308 82 312
rect 36 305 40 308
rect 58 305 62 308
rect 78 305 82 308
rect 36 285 38 305
rect 48 282 52 285
rect 29 278 52 282
rect 48 275 52 278
rect 68 282 72 285
rect 68 278 91 282
rect 68 275 72 278
rect 37 265 38 275
rect 52 265 58 275
rect 78 262 82 265
rect 6 258 43 262
rect 47 258 82 262
rect 67 251 83 255
rect 57 238 58 248
rect 82 238 83 248
rect 42 235 46 236
rect 68 235 72 238
rect 0 231 33 235
rect 37 231 110 235
rect 0 227 110 231
rect 40 220 41 224
rect 58 222 62 227
rect 78 222 80 227
rect 41 211 45 212
rect 48 204 52 212
rect 68 204 72 212
rect 77 204 81 205
rect 38 191 42 194
rect 57 191 60 194
rect 0 187 25 191
rect 38 187 60 191
rect 67 187 110 191
rect 38 184 42 187
rect 57 184 60 187
rect 38 149 42 164
rect 48 152 52 164
rect 61 157 62 161
rect 69 152 72 164
rect 38 145 41 149
rect 39 130 43 131
rect 58 130 62 133
rect 78 130 82 133
rect 0 122 110 130
rect 28 99 32 122
rect 51 114 55 115
rect 58 107 62 122
rect 65 114 69 115
rect 88 107 92 122
rect 28 72 32 86
rect 39 79 43 90
rect 48 79 52 87
rect 68 86 72 87
rect 78 79 82 87
rect 48 75 82 79
rect 68 72 72 75
rect 88 72 92 87
rect 16 52 18 72
rect 82 68 92 72
rect 87 57 91 61
rect 16 42 20 52
rect 58 49 62 52
rect 27 45 62 49
rect 78 45 79 49
rect 58 42 62 45
rect 16 32 18 42
rect 82 32 92 36
rect 16 31 20 32
rect 28 21 32 32
rect 68 29 72 32
rect 39 25 41 29
rect 48 25 82 29
rect 28 4 32 8
rect 48 17 52 25
rect 68 17 72 18
rect 78 17 82 25
rect 88 17 92 32
rect 58 4 62 7
rect 88 4 92 7
rect 0 0 110 4
<< metal2 >>
rect 0 204 6 258
rect 23 216 27 356
rect 36 312 40 336
rect 33 235 37 265
rect 53 248 57 322
rect 83 255 87 322
rect 83 248 87 251
rect 91 233 95 278
rect 69 229 95 233
rect 69 224 73 229
rect 37 220 41 224
rect 45 220 73 224
rect 23 212 41 216
rect 45 212 81 216
rect 77 209 81 212
rect 25 133 29 187
rect 33 157 57 161
rect 33 141 37 157
rect 45 145 67 149
rect 33 137 57 141
rect 25 129 35 133
rect 31 86 35 129
rect 53 119 57 137
rect 55 115 57 119
rect 63 119 67 145
rect 63 115 65 119
rect 43 90 91 94
rect 31 82 68 86
rect 16 0 20 27
rect 41 14 45 25
rect 68 22 72 82
rect 87 65 91 90
rect 79 14 83 45
rect 41 10 83 14
<< ntransistor >>
rect 44 265 46 275
rect 64 265 66 275
rect 74 265 76 275
rect 64 238 66 248
rect 74 238 76 248
rect 54 212 56 222
rect 64 212 66 222
rect 74 212 76 222
rect 44 194 46 204
rect 64 194 66 204
rect 24 32 26 42
rect 34 32 36 42
rect 44 32 46 42
rect 54 32 56 42
rect 64 32 66 42
rect 74 32 76 42
rect 54 7 56 17
rect 64 7 66 17
rect 84 7 86 17
<< ptransistor >>
rect 64 322 66 342
rect 74 322 76 342
rect 44 285 46 305
rect 64 285 66 305
rect 74 285 76 305
rect 44 164 46 184
rect 64 164 66 184
rect 54 133 56 152
rect 64 133 66 152
rect 74 133 76 152
rect 54 87 56 107
rect 64 87 66 107
rect 84 87 86 107
rect 24 52 26 72
rect 34 52 36 72
rect 44 52 46 72
rect 54 52 56 72
rect 64 52 66 72
rect 74 52 76 72
<< polycontact >>
rect 43 308 47 312
rect 73 315 77 319
rect 43 258 47 262
rect 63 251 67 255
rect 36 220 40 224
rect 41 207 45 211
rect 77 200 81 204
rect 63 187 67 191
rect 62 157 66 161
rect 51 110 55 114
rect 65 110 69 114
rect 39 75 43 79
rect 87 53 91 57
rect 23 45 27 49
rect 74 45 78 49
rect 35 25 39 29
<< ndcontact >>
rect 38 265 42 275
rect 48 265 52 275
rect 58 265 62 275
rect 68 265 72 275
rect 78 265 82 275
rect 58 238 62 248
rect 68 238 72 248
rect 78 238 82 248
rect 48 212 52 222
rect 58 212 62 222
rect 68 212 72 222
rect 78 212 82 222
rect 38 194 42 204
rect 48 194 52 204
rect 57 194 62 204
rect 68 194 72 204
rect 18 32 22 42
rect 28 32 32 42
rect 38 32 42 42
rect 48 32 52 42
rect 58 32 62 42
rect 68 32 72 42
rect 78 32 82 42
rect 48 7 52 17
rect 58 7 62 17
rect 68 7 72 17
rect 78 7 82 17
rect 88 7 92 17
<< pdcontact >>
rect 58 322 62 342
rect 68 322 72 342
rect 78 322 82 342
rect 38 285 42 305
rect 48 285 52 305
rect 58 285 62 305
rect 68 285 72 305
rect 78 285 82 305
rect 38 164 42 184
rect 48 164 52 184
rect 57 164 62 184
rect 68 164 72 184
rect 48 133 52 152
rect 58 133 62 152
rect 68 133 72 152
rect 78 133 82 152
rect 48 87 52 107
rect 58 87 62 107
rect 68 87 72 107
rect 78 87 82 107
rect 88 87 92 107
rect 18 52 22 72
rect 28 52 32 72
rect 38 52 42 72
rect 48 52 52 72
rect 58 52 62 72
rect 68 52 72 72
rect 78 52 82 72
<< m2contact >>
rect 36 336 40 340
rect 53 322 57 342
rect 83 322 87 342
rect 36 308 40 312
rect 91 278 95 282
rect 33 265 37 275
rect 0 258 6 262
rect 83 251 87 255
rect 53 238 57 248
rect 83 238 87 248
rect 33 231 37 235
rect 41 220 45 224
rect 41 212 45 216
rect 77 205 81 209
rect 25 187 29 191
rect 57 157 61 161
rect 41 145 45 149
rect 51 115 55 119
rect 65 115 69 119
rect 39 90 43 94
rect 68 82 72 86
rect 87 61 91 65
rect 79 45 83 49
rect 16 27 20 31
rect 41 25 45 29
rect 68 18 72 22
<< psubstratepcontact >>
rect 42 236 46 244
rect 80 222 84 227
rect 28 8 32 21
<< nsubstratencontact >>
rect 43 336 47 344
rect 39 131 43 136
rect 28 86 32 99
<< labels >>
rlabel polysilicon 44 72 46 126 1 BxnorAdd
rlabel metal2 31 82 35 126 1 Cout
rlabel metal2 53 119 57 126 5 Cin
rlabel metal2 63 119 67 126 5 X
rlabel metal2 16 0 20 27 3 sum
rlabel metal2 69 220 73 231 1 BxnorAdd
rlabel metal1 38 187 60 191 1 X
rlabel polysilicon 64 184 66 187 1 Cin
rlabel metal2 91 231 95 278 1 BxnorAdd
rlabel metal1 90 315 94 326 1 AddIn
rlabel metal1 21 187 25 191 3 Cout
rlabel metal2 23 262 27 356 1 A
rlabel metal1 0 322 53 326 1 AddOut
<< end >>
