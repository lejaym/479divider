magic
tech scmos
timestamp 1428729039
<< pwell >>
rect 993 1566 1103 1570
rect 993 1561 1229 1566
rect 993 1548 1653 1561
rect 993 1545 1229 1548
rect 993 1542 1101 1545
rect 1425 1370 1438 1380
rect 902 1185 926 1267
rect 1428 1166 1441 1171
rect 1727 986 1773 1068
<< nwell >>
rect 903 1121 926 1181
rect 909 1116 926 1121
rect 1711 1071 1773 1117
<< polysilicon >>
rect 1707 1433 1715 1434
rect 1710 1329 1712 1433
rect 1730 1410 1732 1434
rect 1740 1410 1742 1434
rect 1730 1328 1732 1365
rect 1740 1329 1742 1362
rect 912 1198 914 1200
rect 912 1178 914 1188
rect 912 1156 914 1158
rect 1754 1097 1755 1101
rect 1735 1093 1737 1095
rect 1753 1093 1755 1097
rect 1763 1097 1764 1101
rect 1763 1093 1765 1097
rect 1735 1072 1737 1075
rect 1735 1068 1736 1072
rect 1735 1065 1737 1068
rect 1753 1065 1755 1075
rect 1763 1065 1765 1075
rect 1735 1053 1737 1055
rect 1753 1053 1755 1055
rect 1763 1053 1765 1055
<< ndiffusion >>
rect 910 1188 912 1198
rect 914 1188 916 1198
rect 1733 1055 1735 1065
rect 1737 1055 1739 1065
rect 1751 1055 1753 1065
rect 1755 1055 1757 1065
rect 1761 1055 1763 1065
rect 1765 1055 1767 1065
<< pdiffusion >>
rect 910 1158 912 1178
rect 914 1158 916 1178
rect 1733 1075 1735 1093
rect 1737 1075 1739 1093
rect 1751 1075 1753 1093
rect 1755 1075 1757 1093
rect 1761 1075 1763 1093
rect 1765 1075 1767 1093
<< metal1 >>
rect 870 2018 1715 2026
rect 870 1888 878 2018
rect 928 2006 1704 2014
rect 20 1880 878 1888
rect 882 1984 998 2000
rect 1645 1984 1689 2000
rect 882 1876 916 1984
rect 1420 1946 1429 1952
rect -36 1840 916 1876
rect 938 1910 1001 1926
rect -35 1778 5 1840
rect 43 1821 49 1828
rect 938 1823 976 1910
rect 910 1807 976 1823
rect -34 1749 4 1778
rect -34 1733 30 1749
rect -34 1560 4 1733
rect 938 1725 976 1807
rect 1665 1799 1689 1984
rect 1642 1783 1689 1799
rect 1424 1742 1430 1751
rect 938 1709 1001 1725
rect 938 1675 976 1709
rect 909 1659 976 1675
rect 915 1635 920 1643
rect 910 1617 917 1623
rect 938 1577 976 1659
rect 1665 1651 1689 1783
rect 1642 1635 1689 1651
rect 938 1561 1000 1577
rect 1096 1561 1229 1566
rect -34 1544 30 1560
rect 938 1554 1653 1561
rect -34 1359 4 1544
rect 938 1538 1002 1554
rect 1096 1545 1229 1554
rect 910 1446 929 1454
rect 938 1433 976 1538
rect 1336 1477 1344 1494
rect 1665 1480 1689 1635
rect 1642 1464 1647 1480
rect 1654 1464 1689 1480
rect 910 1417 976 1433
rect 938 1406 976 1417
rect 1675 1418 1689 1464
rect 1696 1431 1704 2006
rect 1707 1442 1715 2018
rect 1696 1423 1764 1431
rect 1675 1414 1711 1418
rect 938 1390 999 1406
rect 1655 1390 1670 1406
rect 1682 1398 1707 1411
rect -34 1339 30 1359
rect -34 1124 4 1339
rect 938 1229 976 1390
rect 1661 1381 1688 1390
rect 1699 1387 1707 1398
rect 1699 1383 1711 1387
rect 1424 1372 1433 1375
rect 1427 1371 1433 1372
rect 1671 1363 1680 1372
rect 1684 1366 1688 1381
rect 1684 1362 1712 1366
rect 1756 1348 1764 1423
rect 1775 1314 1824 1318
rect 1775 1291 1793 1295
rect 1779 1260 1786 1264
rect 910 1221 976 1229
rect 916 1198 920 1221
rect 938 1205 976 1221
rect 991 1218 999 1226
rect 938 1189 998 1205
rect 1778 1189 1782 1193
rect 906 1178 910 1188
rect 918 1181 921 1185
rect 916 1124 920 1158
rect -34 1116 30 1124
rect 907 1116 920 1124
rect -34 893 4 1116
rect 20 1022 48 1039
rect 938 1021 976 1189
rect 1743 1115 1746 1116
rect 1743 1100 1747 1115
rect 1739 1096 1747 1100
rect 1750 1101 1754 1105
rect 1739 1093 1743 1096
rect 1757 1093 1761 1117
rect 1768 1097 1772 1101
rect 1729 1065 1733 1075
rect 1747 1072 1751 1075
rect 1767 1072 1771 1075
rect 1740 1068 1771 1072
rect 1747 1065 1751 1068
rect 987 1049 1513 1052
rect 1729 1049 1733 1055
rect 987 1044 1733 1049
rect 1739 1044 1743 1055
rect 1767 1044 1771 1055
rect 1739 1040 1771 1044
rect 987 1028 1744 1036
rect 1755 1021 1759 1040
rect 1782 1036 1786 1189
rect 1789 1101 1793 1291
rect 1770 1028 1786 1036
rect 1796 1028 1800 1256
rect 1804 1028 1808 1264
rect 1812 1028 1816 1158
rect 1820 1028 1824 1314
rect 1828 1028 1836 1105
rect 1844 1028 1852 1344
rect 938 998 1865 1021
rect 910 997 1865 998
rect 909 993 1865 997
rect 1785 986 1865 993
rect -34 878 30 893
rect -34 670 4 878
rect 1828 785 1865 986
rect 1787 769 1865 785
rect 1795 745 1796 753
rect 1790 727 1804 733
rect -34 654 30 670
rect -34 524 4 654
rect 1828 555 1865 769
rect 1790 547 1865 555
rect -34 513 30 524
rect -34 385 4 513
rect 1828 459 1865 547
rect 1787 443 1865 459
rect -34 369 30 385
rect -34 237 4 369
rect 1828 311 1865 443
rect 1790 295 1865 311
rect 1790 267 1798 277
rect -34 220 30 237
rect -34 36 4 220
rect 1790 123 1798 131
rect 1828 110 1865 295
rect 1790 94 1865 110
rect -34 20 31 36
rect 1828 19 1865 94
<< metal2 >>
rect 12 1039 20 1880
rect 43 1833 49 1864
rect 43 1823 49 1828
rect 153 1834 159 1864
rect 153 1823 159 1829
rect 263 1833 269 1864
rect 263 1823 269 1828
rect 373 1834 379 1864
rect 373 1823 379 1829
rect 483 1834 489 1864
rect 483 1823 489 1829
rect 593 1833 599 1864
rect 593 1823 599 1828
rect 703 1833 709 1864
rect 703 1823 709 1828
rect 813 1833 819 1864
rect 813 1823 819 1828
rect 920 1643 928 2006
rect 1011 2013 1110 2017
rect 1011 1953 1024 2013
rect 925 1635 928 1643
rect 917 1336 925 1617
rect 1104 1605 1110 2013
rect 1121 2012 1220 2017
rect 1121 1956 1134 2012
rect 1214 1605 1220 2012
rect 1231 2012 1330 2017
rect 1231 1956 1244 2012
rect 1324 1605 1330 2012
rect 1341 2012 1440 2017
rect 1341 1956 1354 2012
rect 1387 1984 1421 1990
rect 1415 1952 1421 1984
rect 1411 1945 1421 1952
rect 1104 1599 1124 1605
rect 1214 1599 1229 1605
rect 1324 1599 1344 1605
rect 995 1565 1011 1571
rect 935 1446 991 1454
rect 917 1328 949 1336
rect 910 1316 933 1320
rect 925 1036 933 1316
rect 941 1052 949 1328
rect 981 1226 991 1446
rect 995 1167 1001 1565
rect 1010 1544 1111 1550
rect 1118 1544 1222 1548
rect 1105 1168 1111 1544
rect 1216 1168 1222 1544
rect 1229 1542 1333 1548
rect 1327 1169 1333 1542
rect 1424 1381 1430 1731
rect 1434 1605 1440 2012
rect 1451 2012 1550 2017
rect 1451 1956 1464 2012
rect 1544 1605 1550 2012
rect 1561 1956 1574 2017
rect 1594 1986 1607 2029
rect 1661 1889 1696 1897
rect 1661 1743 1682 1753
rect 1434 1599 1454 1605
rect 1544 1599 1564 1605
rect 1647 1332 1654 1464
rect 1674 1411 1682 1743
rect 1686 1348 1696 1889
rect 1653 1316 1673 1332
rect 1786 1264 1804 1268
rect 1778 1256 1796 1260
rect 1778 1158 1812 1162
rect 1755 1135 1865 1139
rect 1754 1105 1828 1112
rect 1779 1097 1789 1101
rect 1005 1088 1869 1092
rect 941 1044 979 1052
rect 925 1028 979 1036
rect 1005 994 1011 1088
rect 1115 1080 1869 1084
rect 1115 994 1121 1080
rect 1225 1072 1869 1076
rect 1225 994 1231 1072
rect 1335 1064 1869 1068
rect 1335 994 1341 1064
rect 1445 1056 1869 1060
rect 1445 994 1451 1056
rect 1555 1048 1869 1052
rect 1555 994 1561 1048
rect 1665 1040 1869 1044
rect 1665 994 1671 1040
rect 1752 1028 1762 1036
rect 1774 1032 1869 1036
rect 1774 994 1780 1032
rect 1796 753 1800 1024
rect 1804 733 1808 1024
rect 1812 501 1816 1024
rect 1790 493 1812 501
rect 1820 469 1824 1024
rect 1790 466 1820 469
rect 1794 462 1820 466
rect 1828 277 1836 1024
rect 1806 267 1836 277
rect 1844 131 1852 1024
rect 1804 123 1852 131
rect 81 17 94 20
rect 81 -21 94 11
rect 191 17 204 20
rect 191 -21 204 11
rect 301 17 314 20
rect 301 -21 314 11
rect 411 17 424 20
rect 411 -21 424 11
rect 521 17 534 20
rect 521 -21 534 11
rect 631 17 644 20
rect 631 -21 644 11
rect 741 17 754 20
rect 741 -21 754 11
rect 851 17 864 20
rect 851 -21 864 11
rect 961 17 974 20
rect 961 -21 974 11
rect 1071 17 1084 20
rect 1071 -21 1084 11
rect 1181 17 1194 20
rect 1181 -21 1194 11
rect 1291 17 1304 20
rect 1291 -21 1304 11
rect 1401 17 1414 20
rect 1401 -21 1414 11
rect 1511 17 1524 20
rect 1511 -21 1524 11
rect 1621 17 1634 20
rect 1621 -21 1634 11
rect 1731 17 1744 20
rect 1731 -21 1744 11
<< ntransistor >>
rect 912 1188 914 1198
rect 1735 1055 1737 1065
rect 1753 1055 1755 1065
rect 1763 1055 1765 1065
<< ptransistor >>
rect 912 1158 914 1178
rect 1735 1075 1737 1093
rect 1753 1075 1755 1093
rect 1763 1075 1765 1093
<< polycontact >>
rect 910 1635 915 1643
rect 1707 1434 1715 1442
rect 914 1181 918 1185
rect 1750 1097 1754 1101
rect 1764 1097 1768 1101
rect 1736 1068 1740 1072
rect 1790 745 1795 753
<< ndcontact >>
rect 906 1188 910 1198
rect 916 1188 920 1198
rect 1729 1055 1733 1065
rect 1739 1055 1743 1065
rect 1747 1055 1751 1065
rect 1757 1055 1761 1065
rect 1767 1055 1771 1065
<< pdcontact >>
rect 906 1158 910 1178
rect 916 1158 920 1178
rect 1729 1075 1733 1093
rect 1739 1075 1743 1093
rect 1747 1075 1751 1093
rect 1757 1075 1761 1093
rect 1767 1075 1771 1093
<< m2contact >>
rect 1594 2029 1607 2033
rect 920 2006 928 2014
rect 12 1880 20 1888
rect 43 1828 49 1833
rect 153 1829 159 1834
rect 263 1828 269 1833
rect 373 1829 379 1834
rect 483 1829 489 1834
rect 593 1828 599 1833
rect 703 1828 709 1833
rect 813 1828 819 1833
rect 1651 1889 1661 1897
rect 1651 1743 1661 1753
rect 1424 1731 1430 1742
rect 920 1635 925 1643
rect 917 1617 925 1623
rect 929 1446 935 1454
rect 1647 1464 1654 1480
rect 1658 1425 1662 1429
rect 1666 1425 1670 1429
rect 1674 1398 1682 1411
rect 53 1327 57 1333
rect 163 1326 167 1332
rect 273 1328 277 1334
rect 383 1326 387 1332
rect 493 1326 497 1332
rect 603 1326 607 1332
rect 713 1327 717 1333
rect 823 1326 827 1332
rect 904 1316 910 1320
rect 1424 1375 1430 1381
rect 1640 1316 1653 1332
rect 1782 1264 1786 1268
rect 981 1218 991 1226
rect 1782 1189 1786 1193
rect 921 1181 925 1185
rect 12 1022 20 1039
rect 995 1161 1001 1167
rect 1105 1163 1111 1168
rect 1216 1164 1222 1168
rect 1327 1164 1333 1169
rect 1751 1135 1755 1139
rect 1750 1105 1754 1112
rect 1772 1097 1779 1101
rect 979 1044 987 1052
rect 979 1028 987 1036
rect 1744 1028 1752 1036
rect 1804 1264 1808 1268
rect 1789 1097 1793 1101
rect 1796 1256 1800 1260
rect 1762 1028 1770 1036
rect 1796 1024 1800 1028
rect 1804 1024 1808 1028
rect 1812 1158 1816 1162
rect 1812 1024 1816 1028
rect 1820 1024 1824 1028
rect 1828 1105 1836 1112
rect 1828 1024 1836 1028
rect 1844 1024 1852 1028
rect 156 1004 160 1010
rect 266 1003 270 1009
rect 376 1004 380 1010
rect 486 1003 490 1009
rect 596 1005 600 1011
rect 706 1004 710 1010
rect 816 1004 820 1010
rect 1796 745 1800 753
rect 1804 727 1808 733
rect 87 529 95 535
rect 189 529 197 535
rect 315 529 323 535
rect 417 529 425 535
rect 518 529 526 535
rect 645 529 653 535
rect 746 529 754 535
rect 848 529 856 535
rect 949 529 957 535
rect 1076 529 1084 535
rect 1177 529 1185 535
rect 1279 529 1287 535
rect 1405 529 1413 535
rect 1507 529 1515 535
rect 1622 529 1630 535
rect 1737 529 1745 535
rect 1812 493 1816 501
rect 1790 462 1794 466
rect 1820 462 1824 469
rect 1798 267 1806 277
rect 1798 123 1804 131
rect 81 11 94 17
rect 191 11 204 17
rect 301 11 314 17
rect 411 11 424 17
rect 521 11 534 17
rect 631 11 644 17
rect 741 11 754 17
rect 851 11 864 17
rect 961 11 974 17
rect 1071 11 1084 17
rect 1181 11 1194 17
rect 1291 11 1304 17
rect 1401 11 1414 17
rect 1511 11 1524 17
rect 1621 11 1634 17
rect 1731 11 1744 17
use datapathL  datapathL_0
array 0 7 110 0 0 1803
timestamp 1428729039
transform 1 0 30 0 1 562
box 0 -542 110 1261
use rego  rego_2
timestamp 1428724078
transform 1 0 993 0 -1 1840
box 0 -160 110 279
use rego  rego_3
timestamp 1428724078
transform 1 0 1103 0 -1 1840
box 0 -160 110 279
use rego  rego_5
timestamp 1428724078
transform 1 0 1213 0 -1 1840
box 0 -160 110 279
use rego  rego_6
timestamp 1428724078
transform 1 0 1323 0 -1 1840
box 0 -160 110 279
use rego  rego_7
timestamp 1428724078
transform 1 0 1433 0 -1 1840
box 0 -160 110 279
use rego  rego_8
timestamp 1428724078
transform 1 0 1543 0 -1 1840
box 0 -160 110 279
use rego  rego_4
timestamp 1428724078
transform 1 0 993 0 1 1275
box 0 -160 110 279
use ../cells/rego  rego_9
timestamp 1428724078
transform 1 0 1103 0 1 1275
box 0 -160 110 279
use rego  rego_1
timestamp 1428724078
transform 1 0 1213 0 1 1275
box 0 -160 110 279
use rego  rego_0
timestamp 1428724078
transform 1 0 1323 0 1 1275
box 0 -160 110 279
use and  and_0
timestamp 1427941063
transform 1 0 1736 0 1 1385
box -25 -23 14 33
use smlogic  smlogic_0
timestamp 1428724254
transform 1 0 1304 0 1 1193
box 123 -143 548 366
use datapathS  datapathS_0
array 0 7 110 0 0 974
timestamp 1428724254
transform 1 0 910 0 1 562
box 0 -542 110 432
<< labels >>
rlabel metal2 1790 495 1815 499 0 INBIT
rlabel metal1 -34 20 4 1822 0 Vdd
rlabel metal1 1828 19 1865 1021 0 GND
rlabel space 1594 1974 1607 2004 1 valid
rlabel metal2 920 1643 928 2006 1 clk
rlabel space 1753 1119 1766 1121 1 start
rlabel metal2 1751 1135 1865 1139 1 start
rlabel metal1 1844 1028 1852 1344 1 reset
rlabel space 1594 1974 1607 2033 1 valid
rlabel space 1594 1974 1607 2029 1 valid
rlabel m2contact 1594 2029 1607 2033 5 valid
rlabel space 813 1785 819 1864 1 divisorin_0
rlabel m2contact 813 1828 819 1833 1 divisorin_0
rlabel m2contact 703 1828 709 1833 1 divisorin_1
rlabel m2contact 593 1828 599 1833 1 divisorin_2
rlabel m2contact 483 1829 489 1834 1 divisorin_3
rlabel m2contact 373 1829 379 1834 1 divisorin_4
rlabel m2contact 263 1828 269 1833 1 divisorin_5
rlabel m2contact 153 1829 159 1834 1 divisorin_6
rlabel metal2 1774 1032 1869 1036 1 dividendin_0
rlabel metal2 1665 1040 1869 1044 1 dividendin_1
rlabel metal2 1555 1048 1869 1052 1 dividendin_2
rlabel metal2 1445 1056 1869 1060 1 dividendin_3
rlabel metal2 1335 1064 1869 1068 1 dividendin_4
rlabel metal2 1225 1072 1869 1076 1 dividendin_5
rlabel metal2 1115 1080 1869 1084 1 dividendin_6
rlabel metal2 1005 1088 1869 1092 1 dividendin_7
rlabel space 1731 -21 1744 46 1 quotient_0
rlabel m2contact 1731 11 1744 17 1 quotient_0
rlabel m2contact 1621 11 1634 17 1 quotient_1
rlabel m2contact 1511 11 1524 17 1 quotient_2
rlabel m2contact 1401 11 1414 17 1 quotient_3
rlabel m2contact 1291 11 1304 17 1 quotient_4
rlabel m2contact 1181 11 1194 17 1 quotient_5
rlabel m2contact 1071 11 1084 17 1 quotient_6
rlabel m2contact 961 11 974 17 1 quotient_7
rlabel m2contact 81 11 94 17 1 remainder_6
rlabel m2contact 191 11 204 17 1 remainder_5
rlabel m2contact 301 11 314 17 1 remainder_4
rlabel m2contact 411 11 424 17 1 remainder_3
rlabel m2contact 521 11 534 17 1 remainder_2
rlabel m2contact 631 11 644 17 1 remainder_1
rlabel m2contact 741 11 754 17 1 remainder_0
rlabel space 1740 1329 1742 1370 1 SB1
rlabel polysilicon 1740 1410 1742 1434 1 SB1
rlabel polysilicon 1730 1410 1732 1434 1 SB0
rlabel polysilicon 1707 1433 1715 1434 1 sign
rlabel space 1613 1113 1651 1115 1 SB0_out
rlabel metal2 917 1328 925 1617 1 clkload
rlabel space 1666 1342 1670 1559 1 nextsb1
rlabel m2contact 1666 1425 1670 1429 1 nextsb1
rlabel m2contact 1658 1425 1662 1429 1 nextsb0
rlabel m2contact 816 1004 820 1010 1 sum0
rlabel m2contact 706 1004 710 1010 1 sum1
rlabel m2contact 596 1005 600 1011 1 sum2
rlabel m2contact 486 1003 490 1009 1 sum3
rlabel m2contact 376 1004 380 1010 1 sum4
rlabel space 266 989 270 1021 1 sum5
rlabel space 156 989 160 1021 1 sum6
rlabel m2contact 266 1003 270 1009 1 sum5
rlabel m2contact 156 1004 160 1010 1 sum6
rlabel m2contact 823 1326 827 1332 1 divregout0
rlabel m2contact 713 1327 717 1333 1 divregout1
rlabel m2contact 603 1326 607 1332 1 divregout2
rlabel m2contact 493 1326 497 1332 1 divregout3
rlabel m2contact 383 1326 387 1332 1 divregout4
rlabel m2contact 273 1328 277 1334 1 divregout5
rlabel m2contact 163 1326 167 1332 1 divregout6
rlabel m2contact 53 1327 57 1333 1 divregout7
rlabel m2contact 1737 529 1745 535 1 qmuxout0
rlabel m2contact 1622 529 1630 535 1 qmuxout1
rlabel m2contact 1507 529 1515 535 1 qmuxout2
rlabel m2contact 1405 529 1413 535 1 qmuxout3
rlabel m2contact 1279 529 1287 535 1 qmuxout4
rlabel m2contact 1177 529 1185 535 1 qmuxout5
rlabel m2contact 1076 529 1084 535 1 qmuxout6
rlabel m2contact 949 529 957 535 1 qmuxout7
rlabel m2contact 848 529 856 535 1 rmuxout0
rlabel m2contact 746 529 754 535 1 rmuxout1
rlabel m2contact 645 529 653 535 1 rmuxout2
rlabel m2contact 518 529 526 535 1 rmuxout3
rlabel m2contact 417 529 425 535 1 rmuxout4
rlabel m2contact 315 529 323 535 1 rmuxout5
rlabel m2contact 189 529 197 535 1 rmuxout6
rlabel m2contact 87 529 95 535 1 rmuxout7
rlabel metal1 1775 1314 1812 1318 1 shift
rlabel metal1 1775 1291 1789 1295 1 load
rlabel metal2 1786 1264 1804 1268 1 sel1
rlabel metal1 1796 1024 1800 1252 1 sel0
rlabel space 1776 1189 1782 1193 1 add
rlabel metal2 1778 1158 1812 1162 1 inbit
rlabel m2contact 1782 1189 1786 1193 1 add
<< end >>
