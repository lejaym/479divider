magic
tech scmos
timestamp 1428255215
<< pwell >>
rect 0 237 110 279
rect 0 76 110 155
rect 0 -150 110 -61
<< nwell >>
rect 0 155 110 237
rect 0 -61 110 76
rect 0 -201 110 -150
<< polysilicon >>
rect 22 250 24 252
rect 34 250 37 252
rect 74 250 77 252
rect 87 250 106 252
rect 22 223 24 225
rect 44 223 50 225
rect 46 210 50 223
rect 98 225 106 250
rect 61 223 67 225
rect 87 223 89 225
rect 98 219 99 225
rect 105 219 106 225
rect 46 209 66 210
rect 46 206 72 209
rect 22 184 24 186
rect 74 184 76 186
rect 22 162 24 164
rect 74 162 76 164
rect 11 160 24 162
rect 18 150 24 160
rect 11 148 24 150
rect 54 160 76 162
rect 61 150 76 160
rect 54 148 76 150
rect 22 146 24 148
rect 74 146 76 148
rect 22 134 24 136
rect 74 134 76 136
rect 44 111 46 113
rect 82 111 84 113
rect 44 99 46 101
rect 82 99 84 101
rect 5 91 33 99
rect 44 95 69 99
rect 82 95 110 99
rect 44 91 46 93
rect 26 71 33 91
rect 44 79 46 81
rect 64 80 69 95
rect 82 91 84 93
rect 100 91 110 95
rect 44 78 58 79
rect 44 72 46 78
rect 44 71 58 72
rect 44 69 46 71
rect 67 70 69 80
rect 44 47 46 49
rect 64 45 69 70
rect 82 79 84 81
rect 82 73 92 79
rect 82 69 84 73
rect 82 47 84 49
rect 100 45 105 91
rect 44 42 69 45
rect 82 42 105 45
rect 44 40 46 42
rect 82 40 84 42
rect 44 18 46 20
rect 82 18 84 20
rect 65 -4 67 -2
rect 90 -4 92 -2
rect 15 -40 22 -5
rect 25 -24 27 -22
rect 47 -24 56 -22
rect 15 -42 27 -40
rect 47 -42 49 -40
rect 15 -81 22 -42
rect 51 -63 56 -24
rect 65 -45 67 -43
rect 76 -45 81 -19
rect 90 -26 92 -24
rect 90 -29 105 -26
rect 90 -33 92 -31
rect 65 -52 81 -45
rect 50 -71 56 -63
rect 25 -73 27 -71
rect 37 -73 56 -71
rect 76 -57 81 -52
rect 90 -57 92 -53
rect 76 -67 92 -57
rect 15 -83 25 -81
rect 23 -89 25 -83
rect 23 -91 27 -89
rect 37 -91 40 -89
rect 76 -90 81 -67
rect 90 -69 92 -67
rect 90 -81 92 -79
rect 100 -83 105 -29
rect 90 -87 105 -83
rect 90 -89 92 -87
rect 100 -90 105 -87
rect 90 -101 92 -99
rect 33 -131 35 -129
rect 75 -131 77 -129
rect 33 -143 35 -141
rect 75 -143 77 -141
rect 33 -145 50 -143
rect 33 -155 43 -145
rect 33 -157 50 -155
rect 75 -145 88 -143
rect 75 -155 81 -145
rect 75 -157 88 -155
rect 33 -159 35 -157
rect 75 -159 77 -157
rect 33 -181 35 -179
rect 75 -181 77 -179
<< ndiffusion >>
rect 24 252 34 253
rect 24 249 34 250
rect 77 252 87 253
rect 77 249 87 250
rect 21 136 22 146
rect 24 136 25 146
rect 73 136 74 146
rect 76 136 77 146
rect 43 101 44 111
rect 46 101 47 111
rect 81 101 82 111
rect 84 101 85 111
rect 43 81 44 91
rect 46 81 47 91
rect 81 81 82 91
rect 84 81 85 91
rect 27 -71 37 -70
rect 27 -74 37 -73
rect 27 -89 37 -88
rect 89 -79 90 -69
rect 92 -79 93 -69
rect 27 -92 37 -91
rect 89 -99 90 -89
rect 92 -99 93 -89
rect 32 -141 33 -131
rect 35 -141 36 -131
rect 74 -141 75 -131
rect 77 -141 78 -131
<< pdiffusion >>
rect 24 225 44 226
rect 24 222 44 223
rect 67 225 87 226
rect 67 222 87 223
rect 21 164 22 184
rect 24 164 25 184
rect 73 164 74 184
rect 76 164 77 184
rect 43 49 44 69
rect 46 49 47 69
rect 81 49 82 69
rect 84 49 85 69
rect 43 20 44 40
rect 46 20 47 40
rect 81 20 82 40
rect 84 20 85 40
rect 27 -22 47 -21
rect 27 -25 47 -24
rect 27 -40 47 -39
rect 27 -43 47 -42
rect 64 -43 65 -4
rect 67 -43 68 -4
rect 89 -24 90 -4
rect 92 -24 93 -4
rect 89 -53 90 -33
rect 92 -53 93 -33
rect 32 -179 33 -159
rect 35 -179 36 -159
rect 74 -179 75 -159
rect 77 -179 78 -159
<< metal1 >>
rect 0 277 110 279
rect 0 265 14 277
rect 21 265 42 277
rect 49 265 71 277
rect 78 265 110 277
rect 0 263 110 265
rect 10 253 24 257
rect 37 256 53 257
rect 37 255 46 256
rect 10 242 21 253
rect 43 250 46 255
rect 52 250 53 256
rect 87 253 100 257
rect 43 249 53 250
rect 10 235 13 242
rect 20 235 21 242
rect 10 222 21 235
rect 24 241 87 245
rect 24 235 28 241
rect 34 235 87 241
rect 24 230 87 235
rect 10 218 24 222
rect 52 221 55 227
rect 90 240 100 253
rect 96 234 100 240
rect 90 229 100 234
rect 90 222 96 229
rect 52 219 61 221
rect 58 213 61 219
rect 87 218 96 222
rect 105 219 106 225
rect 99 216 106 219
rect 52 212 61 213
rect 72 209 75 215
rect 99 210 100 216
rect 66 208 81 209
rect 0 203 110 205
rect 0 191 16 203
rect 23 191 41 203
rect 48 191 79 203
rect 86 191 110 203
rect 0 189 110 191
rect 13 184 21 189
rect 65 184 73 189
rect 13 164 17 184
rect 29 164 49 184
rect 65 164 69 184
rect 81 164 98 184
rect 37 162 49 164
rect 37 160 61 162
rect 18 158 33 160
rect 18 152 27 158
rect 18 150 33 152
rect 37 150 54 160
rect 37 148 61 150
rect 86 159 98 164
rect 86 153 87 159
rect 93 153 98 159
rect 37 146 49 148
rect 86 146 98 153
rect 13 136 17 146
rect 29 145 49 146
rect 29 138 33 145
rect 40 138 49 145
rect 29 136 49 138
rect 65 136 69 146
rect 81 136 98 146
rect 13 131 21 136
rect 65 131 73 136
rect 0 129 110 131
rect 0 117 14 129
rect 21 117 42 129
rect 49 117 71 129
rect 78 117 110 129
rect 0 115 110 117
rect 47 111 51 115
rect 85 111 89 115
rect 15 109 39 111
rect 15 103 30 109
rect 36 103 39 109
rect 15 101 39 103
rect 15 79 25 101
rect 47 91 51 101
rect 5 73 25 79
rect 15 40 25 73
rect 29 79 39 91
rect 54 101 77 111
rect 29 71 33 79
rect 54 78 60 101
rect 85 91 89 101
rect 58 72 60 78
rect 29 58 39 71
rect 35 52 39 58
rect 29 49 39 52
rect 47 40 51 49
rect 15 20 39 40
rect 54 40 60 72
rect 63 80 81 81
rect 67 77 81 80
rect 67 71 72 77
rect 78 71 81 77
rect 97 73 110 79
rect 67 70 81 71
rect 63 69 81 70
rect 85 40 89 49
rect 54 32 77 40
rect 54 26 57 32
rect 63 26 77 32
rect 54 20 77 26
rect 47 16 51 20
rect 85 16 89 20
rect 0 14 110 16
rect 0 3 16 14
rect 23 3 41 14
rect 48 3 79 14
rect 86 3 110 14
rect 0 0 110 3
rect 68 -4 72 0
rect 93 -4 97 0
rect 30 -11 34 -5
rect 10 -21 27 -17
rect 10 -77 16 -21
rect 47 -29 60 -25
rect 27 -35 60 -29
rect 47 -39 60 -35
rect 22 -47 27 -43
rect 22 -54 37 -47
rect 22 -61 28 -54
rect 35 -61 37 -54
rect 22 -66 37 -61
rect 22 -70 27 -66
rect 48 -57 50 -51
rect 42 -63 50 -57
rect 42 -71 45 -63
rect 53 -56 60 -39
rect 76 -8 85 -4
rect 81 -19 85 -8
rect 76 -24 85 -19
rect 93 -33 97 -24
rect 53 -63 72 -56
rect 53 -69 66 -63
rect 10 -82 22 -77
rect 14 -90 22 -82
rect 53 -78 60 -69
rect 80 -75 85 -33
rect 27 -84 60 -78
rect 64 -84 85 -75
rect 0 -98 11 -90
rect 20 -92 22 -90
rect 20 -96 27 -92
rect 5 -100 11 -98
rect 64 -100 72 -84
rect 93 -89 97 -79
rect 76 -90 85 -89
rect 81 -98 85 -90
rect 76 -99 85 -98
rect 106 -98 110 -90
rect 5 -108 72 -100
rect 93 -111 97 -99
rect 0 -113 110 -111
rect 0 -125 14 -113
rect 21 -125 42 -113
rect 49 -125 71 -113
rect 78 -125 110 -113
rect 0 -127 110 -125
rect 36 -131 44 -127
rect 78 -131 86 -127
rect 11 -141 28 -131
rect 40 -141 44 -131
rect 50 -141 70 -131
rect 82 -141 86 -131
rect 11 -148 23 -141
rect 11 -154 16 -148
rect 22 -154 23 -148
rect 11 -159 23 -154
rect 50 -159 62 -141
rect 66 -147 81 -145
rect 72 -153 81 -147
rect 66 -155 81 -153
rect 11 -179 28 -159
rect 40 -179 44 -159
rect 50 -168 70 -159
rect 50 -175 54 -168
rect 61 -175 70 -168
rect 50 -179 70 -175
rect 82 -179 86 -159
rect 36 -185 44 -179
rect 78 -185 86 -179
rect 0 -187 110 -185
rect 0 -199 16 -187
rect 23 -199 41 -187
rect 48 -199 79 -187
rect 86 -199 110 -187
rect 0 -201 110 -199
<< metal2 >>
rect 12 242 21 279
rect 40 256 53 257
rect 40 250 46 256
rect 52 250 53 256
rect 40 249 53 250
rect 12 235 13 242
rect 20 235 21 242
rect 12 233 21 235
rect 25 241 36 242
rect 25 235 28 241
rect 34 235 36 241
rect 25 158 36 235
rect 40 175 48 249
rect 85 234 90 240
rect 58 213 59 219
rect 52 185 59 213
rect 69 209 75 215
rect 69 206 81 209
rect 52 180 64 185
rect 40 163 53 175
rect 25 152 27 158
rect 33 152 36 158
rect 25 151 36 152
rect 18 145 40 147
rect 18 138 33 145
rect 18 136 40 138
rect 18 -52 25 136
rect 45 111 53 163
rect 30 109 53 111
rect 36 103 53 109
rect 30 101 53 103
rect 57 97 64 180
rect 32 90 64 97
rect 32 58 41 90
rect 69 78 76 206
rect 85 159 96 234
rect 85 153 87 159
rect 93 153 96 159
rect 85 151 96 153
rect 106 210 108 216
rect 69 77 79 78
rect 69 71 72 77
rect 78 71 79 77
rect 69 70 79 71
rect 35 52 41 58
rect 32 -5 41 52
rect 100 34 108 210
rect 32 -11 34 -5
rect 40 -11 41 -5
rect 32 -13 41 -11
rect 55 32 108 34
rect 55 26 57 32
rect 63 26 108 32
rect 55 24 108 26
rect 55 -49 65 24
rect 41 -51 65 -49
rect 18 -54 37 -52
rect 18 -61 28 -54
rect 35 -61 37 -54
rect 41 -57 42 -51
rect 48 -57 65 -51
rect 41 -58 65 -57
rect 18 -63 37 -61
rect 64 -69 66 -63
rect 72 -69 74 -63
rect 20 -96 25 -90
rect 16 -148 25 -96
rect 22 -154 25 -148
rect 64 -147 74 -69
rect 64 -153 66 -147
rect 72 -153 74 -147
rect 64 -154 74 -153
rect 51 -168 64 -165
rect 51 -175 54 -168
rect 61 -175 64 -168
rect 51 -201 64 -175
<< ntransistor >>
rect 24 250 34 252
rect 77 250 87 252
rect 22 136 24 146
rect 74 136 76 146
rect 44 101 46 111
rect 82 101 84 111
rect 44 81 46 91
rect 82 81 84 91
rect 27 -73 37 -71
rect 27 -91 37 -89
rect 90 -79 92 -69
rect 90 -99 92 -89
rect 33 -141 35 -131
rect 75 -141 77 -131
<< ptransistor >>
rect 24 223 44 225
rect 67 223 87 225
rect 22 164 24 184
rect 74 164 76 184
rect 44 49 46 69
rect 82 49 84 69
rect 44 20 46 40
rect 82 20 84 40
rect 27 -24 47 -22
rect 27 -42 47 -40
rect 65 -43 67 -4
rect 90 -24 92 -4
rect 90 -53 92 -33
rect 33 -179 35 -159
rect 75 -179 77 -159
<< polycontact >>
rect 37 249 43 255
rect 55 221 61 227
rect 99 219 105 225
rect 66 209 72 215
rect 11 150 18 160
rect 54 150 61 160
rect 33 71 39 79
rect 46 72 58 78
rect 63 70 67 80
rect 92 73 97 79
rect 22 -11 30 -5
rect 76 -19 81 -8
rect 45 -71 50 -63
rect 76 -98 81 -90
rect 100 -98 106 -90
rect 43 -155 50 -145
rect 81 -155 88 -145
<< ndcontact >>
rect 24 253 34 257
rect 77 253 87 257
rect 24 245 34 249
rect 77 245 87 249
rect 17 136 21 146
rect 25 136 29 146
rect 69 136 73 146
rect 77 136 81 146
rect 39 101 43 111
rect 47 101 51 111
rect 77 101 81 111
rect 85 101 89 111
rect 39 81 43 91
rect 47 81 51 91
rect 77 81 81 91
rect 85 81 89 91
rect 27 -70 37 -66
rect 27 -78 37 -74
rect 27 -88 37 -84
rect 85 -79 89 -69
rect 93 -79 97 -69
rect 27 -96 37 -92
rect 85 -99 89 -89
rect 93 -99 97 -89
rect 28 -141 32 -131
rect 36 -141 40 -131
rect 70 -141 74 -131
rect 78 -141 82 -131
<< pdcontact >>
rect 24 226 44 230
rect 24 218 44 222
rect 67 226 87 230
rect 67 218 87 222
rect 17 164 21 184
rect 25 164 29 184
rect 69 164 73 184
rect 77 164 81 184
rect 39 49 43 69
rect 47 49 51 69
rect 77 49 81 69
rect 85 49 89 69
rect 39 20 43 40
rect 47 20 51 40
rect 77 20 81 40
rect 85 20 89 40
rect 27 -21 47 -17
rect 27 -29 47 -25
rect 27 -39 47 -35
rect 27 -47 47 -43
rect 60 -43 64 -4
rect 68 -43 72 -4
rect 85 -24 89 -4
rect 93 -24 97 -4
rect 85 -53 89 -33
rect 93 -53 97 -33
rect 28 -179 32 -159
rect 36 -179 40 -159
rect 70 -179 74 -159
rect 78 -179 82 -159
<< m2contact >>
rect 46 250 52 256
rect 13 235 20 242
rect 28 235 34 241
rect 90 234 96 240
rect 52 213 58 219
rect 75 209 81 215
rect 100 210 106 216
rect 27 152 33 158
rect 87 153 93 159
rect 33 138 40 145
rect 30 103 36 109
rect 29 52 35 58
rect 72 71 78 77
rect 57 26 63 32
rect 34 -11 40 -5
rect 28 -61 35 -54
rect 42 -57 48 -51
rect 66 -69 72 -63
rect 14 -96 20 -90
rect 16 -154 22 -148
rect 66 -153 72 -147
rect 54 -175 61 -168
<< psubstratepcontact >>
rect 14 265 21 277
rect 42 265 49 277
rect 71 265 78 277
rect 14 117 21 129
rect 42 117 49 129
rect 71 117 78 129
rect 14 -125 21 -113
rect 42 -125 49 -113
rect 71 -125 78 -113
<< nsubstratencontact >>
rect 16 191 23 203
rect 41 191 48 203
rect 79 191 86 203
rect 16 3 23 14
rect 41 3 48 14
rect 79 3 86 14
rect 16 -199 23 -187
rect 41 -199 48 -187
rect 79 -199 86 -187
<< labels >>
rlabel polysilicon 100 -87 105 -67 0 RST
rlabel metal2 51 -201 64 -175 0 REGOUT
rlabel polysilicon 5 91 33 99 0 INCLK
rlabel metal1 5 73 25 79 0 INCLKCLD
rlabel metal2 12 233 21 279 0 REGIN
rlabel polysilicon 100 91 110 99 0 CLK
rlabel metal1 97 73 110 79 0 CLKLD
rlabel metal1 54 32 77 40 0 INCLKn
rlabel polysilicon 64 42 69 70 0 INCLKLDn
rlabel metal1 27 -84 60 -78 0 REGOUTn
rlabel metal1 37 148 54 162 0 REGMEM
<< end >>
