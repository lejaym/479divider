magic
tech scmos
timestamp 1428357410
<< pwell >>
rect -20 399 90 447
rect -20 187 90 280
rect -20 0 90 48
<< nwell >>
rect -20 288 90 391
rect -20 56 90 179
<< polysilicon >>
rect 43 428 64 430
rect 74 428 76 430
rect -4 417 -2 419
rect 6 416 28 418
rect 38 416 40 418
rect -4 404 -2 407
rect -4 398 2 404
rect -1 384 2 398
rect 6 397 10 416
rect 14 410 28 412
rect 38 410 40 412
rect -4 381 2 384
rect -4 378 -2 381
rect -4 356 -2 358
rect 6 355 10 391
rect 14 373 17 410
rect 43 393 49 428
rect 52 412 58 419
rect 52 410 64 412
rect 74 410 76 412
rect 52 401 58 410
rect 52 395 74 401
rect 43 373 49 387
rect 69 388 74 395
rect 69 382 85 388
rect 14 371 19 373
rect 39 371 41 373
rect 43 371 54 373
rect 74 371 76 373
rect 43 355 49 371
rect 79 362 85 382
rect 6 353 19 355
rect 39 353 41 355
rect 43 353 54 355
rect 74 353 76 355
rect 6 322 19 324
rect 39 322 41 324
rect 43 322 54 324
rect 74 322 76 324
rect -4 319 -2 321
rect -4 296 -2 299
rect -4 293 2 296
rect -1 279 2 293
rect 6 286 10 322
rect 43 306 49 322
rect 14 304 19 306
rect 39 304 41 306
rect 43 304 54 306
rect 74 304 76 306
rect -4 273 2 279
rect -4 270 -2 273
rect 6 261 10 280
rect 14 267 17 304
rect 43 290 49 304
rect 79 295 85 315
rect 14 265 28 267
rect 38 265 40 267
rect -4 258 -2 260
rect 6 259 28 261
rect 38 259 40 261
rect 43 249 49 284
rect 52 289 85 295
rect 52 267 58 289
rect 52 265 64 267
rect 74 265 76 267
rect 52 258 58 265
rect 43 247 64 249
rect 74 247 76 249
rect 19 218 21 220
rect 47 218 49 220
rect 19 206 21 208
rect 47 206 49 208
rect -20 198 8 206
rect 19 202 41 206
rect 47 202 90 206
rect 19 198 21 200
rect 1 186 8 198
rect 36 188 41 202
rect 47 198 49 200
rect 65 198 90 202
rect 19 186 21 188
rect 1 185 33 186
rect 1 179 21 185
rect 1 178 33 179
rect 19 176 21 178
rect 40 176 41 188
rect 47 186 49 188
rect 47 180 57 186
rect 47 176 49 180
rect 19 154 21 156
rect 36 152 41 176
rect 47 154 49 156
rect 65 152 70 198
rect 19 149 41 152
rect 47 149 70 152
rect 19 147 21 149
rect 47 147 49 149
rect 19 125 21 127
rect 47 125 49 127
rect -6 92 8 94
rect 28 92 30 94
rect 33 92 43 94
rect 63 92 65 94
rect -6 31 -2 92
rect 33 76 38 92
rect 2 74 8 76
rect 28 74 30 76
rect 33 74 43 76
rect 63 74 65 76
rect 2 37 6 74
rect 33 60 38 74
rect 68 66 74 85
rect 2 35 17 37
rect 27 35 29 37
rect -6 29 17 31
rect 27 29 29 31
rect 33 19 38 54
rect 42 60 74 66
rect 42 37 48 60
rect 42 35 53 37
rect 63 35 65 37
rect 42 28 48 35
rect 33 17 53 19
rect 63 17 65 19
<< ndiffusion >>
rect 64 430 74 431
rect 28 418 38 419
rect -5 407 -4 417
rect -2 407 -1 417
rect 28 412 38 416
rect 28 409 38 410
rect 64 427 74 428
rect 64 412 74 413
rect 64 409 74 410
rect -5 260 -4 270
rect -2 260 -1 270
rect 28 267 38 268
rect 28 261 38 265
rect 28 258 38 259
rect 64 267 74 268
rect 64 264 74 265
rect 64 249 74 250
rect 64 246 74 247
rect 18 208 19 218
rect 21 208 22 218
rect 46 208 47 218
rect 49 208 50 218
rect 18 188 19 198
rect 21 188 22 198
rect 46 188 47 198
rect 49 188 50 198
rect 17 37 27 38
rect 17 31 27 35
rect 17 28 27 29
rect 53 37 63 38
rect 53 34 63 35
rect 53 19 63 20
rect 53 16 63 17
<< pdiffusion >>
rect -5 358 -4 378
rect -2 358 -1 378
rect 19 373 39 374
rect 54 373 74 374
rect 19 370 39 371
rect 19 355 39 356
rect 54 370 74 371
rect 54 355 74 356
rect 19 352 39 353
rect 54 352 74 353
rect 19 324 39 325
rect 54 324 74 325
rect -5 299 -4 319
rect -2 299 -1 319
rect 19 321 39 322
rect 19 306 39 307
rect 54 321 74 322
rect 54 306 74 307
rect 19 303 39 304
rect 54 303 74 304
rect 18 156 19 176
rect 21 156 22 176
rect 46 156 47 176
rect 49 156 50 176
rect 18 127 19 147
rect 21 127 22 147
rect 46 127 47 147
rect 49 127 50 147
rect 8 94 28 95
rect 43 94 63 95
rect 8 91 28 92
rect 8 76 28 77
rect 43 91 63 92
rect 43 76 63 77
rect 8 73 28 74
rect 43 73 63 74
<< metal1 >>
rect -20 445 90 447
rect -20 441 8 445
rect 15 441 29 445
rect 36 441 51 445
rect 58 441 90 445
rect -20 439 90 441
rect -10 417 -5 439
rect 28 423 38 439
rect 64 435 74 439
rect 58 423 64 425
rect 58 420 74 423
rect -10 407 -9 417
rect 3 407 11 417
rect 74 413 85 417
rect -10 392 -4 398
rect 5 397 11 407
rect 19 391 25 396
rect 5 385 11 391
rect 23 385 25 391
rect 28 393 38 405
rect 54 405 64 409
rect 28 387 43 393
rect 28 385 49 387
rect -1 381 11 385
rect -1 378 3 381
rect 10 374 19 378
rect -9 346 -5 358
rect 10 352 16 374
rect 43 366 49 385
rect 54 391 74 405
rect 78 399 85 413
rect 54 383 58 391
rect 66 383 74 391
rect 54 378 74 383
rect 78 370 85 391
rect 74 366 85 370
rect 19 360 49 366
rect 74 356 79 360
rect 10 348 19 352
rect 10 346 39 348
rect 54 346 74 348
rect -20 344 90 346
rect -20 333 -3 344
rect 4 333 22 344
rect 29 333 60 344
rect 67 333 90 344
rect -20 331 90 333
rect -9 319 -5 331
rect 10 329 39 331
rect 10 325 19 329
rect 54 329 74 331
rect 10 303 16 325
rect 74 317 79 321
rect 19 311 49 317
rect 10 299 19 303
rect -1 296 3 299
rect -1 292 11 296
rect 43 292 49 311
rect 74 307 85 311
rect -10 279 -4 285
rect 5 286 11 292
rect 23 286 25 292
rect 5 270 11 280
rect 19 281 25 286
rect 28 290 49 292
rect 28 284 43 290
rect 54 286 74 299
rect 78 286 85 307
rect -10 260 -9 270
rect 3 260 11 270
rect 28 272 38 284
rect 54 278 64 286
rect 72 278 74 286
rect 54 272 74 278
rect 54 268 64 272
rect 78 264 85 278
rect 74 260 85 264
rect -10 238 -5 260
rect 28 238 38 254
rect 58 254 74 257
rect 58 252 64 254
rect 64 238 74 242
rect -20 236 90 238
rect -20 224 -6 236
rect 1 224 22 236
rect 29 224 51 236
rect 58 224 90 236
rect -20 222 90 224
rect 22 218 26 222
rect 50 218 54 222
rect -10 208 14 218
rect -10 186 0 208
rect 22 198 26 208
rect -20 180 0 186
rect -10 147 0 180
rect 4 185 14 198
rect 29 208 42 218
rect 29 185 33 208
rect 50 198 54 208
rect 38 188 42 198
rect 4 179 9 185
rect 4 156 14 179
rect 22 147 26 156
rect -10 137 14 147
rect -10 131 -2 137
rect 4 131 14 137
rect -10 127 14 131
rect 29 147 33 179
rect 40 176 42 188
rect 62 180 90 186
rect 38 156 42 176
rect 50 147 54 156
rect 29 127 42 147
rect 22 123 26 127
rect 50 123 54 127
rect -20 121 90 123
rect -20 110 -4 121
rect 3 110 21 121
rect 28 110 59 121
rect 66 110 90 121
rect -20 107 90 110
rect -3 99 3 107
rect 43 99 63 107
rect -3 95 8 99
rect -3 73 3 95
rect 63 87 68 91
rect 8 81 38 87
rect -3 69 8 73
rect 32 64 38 81
rect 63 77 81 81
rect 8 51 14 56
rect 12 45 14 51
rect 17 60 38 64
rect 17 54 32 60
rect 17 42 27 54
rect 30 44 38 54
rect 43 57 63 69
rect 43 49 52 57
rect 60 49 63 57
rect 43 42 63 49
rect 43 38 53 42
rect 68 50 81 77
rect 68 42 72 50
rect 80 42 81 50
rect 68 34 81 42
rect 63 30 81 34
rect -6 17 0 23
rect 17 8 27 24
rect 48 24 63 27
rect 48 22 53 24
rect 53 8 63 12
rect -20 6 90 8
rect -20 2 8 6
rect 15 2 45 6
rect 52 2 66 6
rect 73 2 90 6
rect -20 0 90 2
<< metal2 >>
rect -10 407 40 415
rect -10 392 -2 407
rect -4 386 -2 392
rect 16 396 19 402
rect 25 396 26 402
rect 16 368 26 396
rect -4 359 26 368
rect -4 294 4 359
rect 32 339 40 407
rect -10 291 4 294
rect -4 285 4 291
rect -10 283 4 285
rect -4 137 4 283
rect -4 131 -2 137
rect -4 20 4 131
rect 9 332 40 339
rect 9 283 17 332
rect 45 286 53 447
rect 58 441 81 447
rect 58 391 66 441
rect 76 391 77 399
rect 76 286 85 391
rect 9 281 25 283
rect 9 275 19 281
rect 45 278 64 286
rect 76 278 77 286
rect 9 273 25 275
rect 9 185 17 273
rect 15 179 17 185
rect 9 62 17 179
rect 14 56 17 62
rect 8 55 17 56
rect -6 17 4 20
rect 0 11 4 17
rect 37 49 52 57
rect 76 50 85 278
rect 37 0 45 49
rect 80 42 85 50
rect 76 0 85 42
<< ntransistor >>
rect 64 428 74 430
rect -4 407 -2 417
rect 28 416 38 418
rect 28 410 38 412
rect 64 410 74 412
rect -4 260 -2 270
rect 28 265 38 267
rect 28 259 38 261
rect 64 265 74 267
rect 64 247 74 249
rect 19 208 21 218
rect 47 208 49 218
rect 19 188 21 198
rect 47 188 49 198
rect 17 35 27 37
rect 17 29 27 31
rect 53 35 63 37
rect 53 17 63 19
<< ptransistor >>
rect -4 358 -2 378
rect 19 371 39 373
rect 54 371 74 373
rect 19 353 39 355
rect 54 353 74 355
rect 19 322 39 324
rect 54 322 74 324
rect -4 299 -2 319
rect 19 304 39 306
rect 54 304 74 306
rect 19 156 21 176
rect 47 156 49 176
rect 19 127 21 147
rect 47 127 49 147
rect 8 92 28 94
rect 43 92 63 94
rect 8 74 28 76
rect 43 74 63 76
<< polycontact >>
rect -10 398 -4 404
rect 5 391 11 397
rect 52 419 58 425
rect 17 385 23 391
rect 43 387 49 393
rect 79 356 85 362
rect 79 315 85 321
rect 5 280 11 286
rect -10 273 -4 279
rect 17 286 23 292
rect 43 284 49 290
rect 52 252 58 258
rect 21 179 33 185
rect 36 176 40 188
rect 57 180 62 186
rect 68 85 74 91
rect 32 54 38 60
rect 6 45 12 51
rect -6 23 0 29
rect 42 22 48 28
<< ndcontact >>
rect 64 431 74 435
rect 28 419 38 423
rect -9 407 -5 417
rect -1 407 3 417
rect 28 405 38 409
rect 64 423 74 427
rect 64 413 74 417
rect 64 405 74 409
rect -9 260 -5 270
rect -1 260 3 270
rect 28 268 38 272
rect 28 254 38 258
rect 64 268 74 272
rect 64 260 74 264
rect 64 250 74 254
rect 64 242 74 246
rect 14 208 18 218
rect 22 208 26 218
rect 42 208 46 218
rect 50 208 54 218
rect 14 188 18 198
rect 22 188 26 198
rect 42 188 46 198
rect 50 188 54 198
rect 17 38 27 42
rect 17 24 27 28
rect 53 38 63 42
rect 53 30 63 34
rect 53 20 63 24
rect 53 12 63 16
<< pdcontact >>
rect -9 358 -5 378
rect -1 358 3 378
rect 19 374 39 378
rect 54 374 74 378
rect 19 366 39 370
rect 19 356 39 360
rect 54 366 74 370
rect 54 356 74 360
rect 19 348 39 352
rect 54 348 74 352
rect 19 325 39 329
rect 54 325 74 329
rect -9 299 -5 319
rect -1 299 3 319
rect 19 317 39 321
rect 19 307 39 311
rect 54 317 74 321
rect 54 307 74 311
rect 19 299 39 303
rect 54 299 74 303
rect 14 156 18 176
rect 22 156 26 176
rect 42 156 46 176
rect 50 156 54 176
rect 14 127 18 147
rect 22 127 26 147
rect 42 127 46 147
rect 50 127 54 147
rect 8 95 28 99
rect 43 95 63 99
rect 8 87 28 91
rect 8 77 28 81
rect 43 87 63 91
rect 43 77 63 81
rect 8 69 28 73
rect 43 69 63 73
<< m2contact >>
rect -10 386 -4 392
rect 19 396 25 402
rect 77 391 85 399
rect 58 383 66 391
rect -10 285 -4 291
rect 19 275 25 281
rect 64 278 72 286
rect 77 278 85 286
rect 9 179 15 185
rect -2 131 4 137
rect 8 56 14 62
rect 52 49 60 57
rect 72 42 80 50
rect -6 11 0 17
<< psubstratepcontact >>
rect 8 441 15 445
rect 29 441 36 445
rect 51 441 58 445
rect -6 224 1 236
rect 22 224 29 236
rect 51 224 58 236
rect 8 2 15 6
rect 45 2 52 6
rect 66 2 73 6
<< nsubstratencontact >>
rect -3 333 4 344
rect 22 333 29 344
rect 60 333 67 344
rect -4 110 3 121
rect 21 110 28 121
rect 59 110 66 121
<< labels >>
rlabel metal1 62 181 77 185 0 S1
rlabel polysilicon 70 198 85 206 0 S0
rlabel metal2 76 115 85 345 0 MUXOUT
rlabel metal2 37 0 45 57 0 REGIN
rlabel metal2 76 50 85 278 0 MUXOUT
rlabel m2contact 64 278 72 286 0 ADDSUB
rlabel metal1 -15 0 8 8 0 GND
rlabel metal1 28 107 59 123 0 Vdd
rlabel m2contact 58 383 66 391 0 DIVIN
<< end >>
