magic
tech scmos
timestamp 1428724254
<< pwell >>
rect 0 690 38 700
rect 6 684 38 690
rect 17 676 38 684
<< metal2 >>
rect 27 781 54 788
rect 0 -15 6 670
rect 16 427 65 432
rect 0 -21 65 -15
rect 4 -493 10 -21
rect 96 -27 105 -15
rect 27 -33 105 -27
rect 27 -45 31 -33
rect 37 -105 41 -103
rect 21 -110 41 -105
rect 4 -500 31 -493
<< m2contact >>
rect 95 426 101 432
use reg  reg_0 ../cells
timestamp 1428354897
transform 1 0 18 0 1 982
box -18 -201 92 279
use adder  adder_0 ../cells
timestamp 1428713239
transform 1 0 0 0 1 432
box 0 0 110 356
use mux  mux_0 ../cells
timestamp 1428357410
transform 1 0 20 0 1 -15
box -20 0 90 447
use shifter  shifter_0 ../cells
timestamp 1428356401
transform 1 0 35 0 1 -106
box -35 3 75 68
use rego  rego_0 ../cells
timestamp 1428724078
transform 1 0 0 0 1 -382
box 0 -160 110 279
<< end >>
