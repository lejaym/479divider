magic
tech scmos
timestamp 1428629792
<< pwell >>
rect 903 1221 910 1234
rect 900 1185 939 1214
<< nwell >>
rect 908 1153 940 1181
rect 903 1124 940 1153
<< polysilicon >>
rect 912 1199 918 1201
rect 928 1199 944 1201
rect 940 1184 944 1199
rect 940 1178 942 1184
rect 940 1157 944 1178
rect 915 1155 917 1157
rect 935 1155 946 1157
<< ndiffusion >>
rect 918 1201 928 1203
rect 918 1197 928 1199
<< pdiffusion >>
rect 917 1157 935 1159
rect 917 1153 935 1155
<< metal1 >>
rect 49 1856 116 1864
rect 159 1859 226 1867
rect 269 1856 336 1864
rect 379 1856 446 1864
rect 489 1856 556 1864
rect 599 1856 666 1864
rect 709 1856 776 1864
rect 819 1856 886 1864
rect -34 1749 4 1822
rect 910 1807 976 1823
rect -34 1733 30 1749
rect -34 1560 4 1733
rect 938 1675 976 1807
rect 909 1659 976 1675
rect 915 1635 920 1643
rect 910 1617 920 1623
rect -34 1544 30 1560
rect -34 1359 4 1544
rect 910 1446 919 1454
rect 938 1433 976 1659
rect 910 1417 976 1433
rect -34 1339 30 1359
rect -34 1124 4 1339
rect 938 1262 976 1417
rect 1912 1424 1936 1484
rect 938 1229 1003 1262
rect 910 1221 1003 1229
rect 918 1209 928 1221
rect 938 1218 1003 1221
rect 910 1166 928 1191
rect 948 1178 956 1190
rect 903 1124 917 1153
rect -34 1116 30 1124
rect 966 1123 1004 1218
rect -34 893 4 1116
rect 938 1092 1000 1123
rect 938 1021 976 1092
rect 1012 1064 1079 1072
rect 1123 1064 1190 1072
rect 1233 1063 1300 1071
rect 1343 1066 1410 1074
rect 1454 1065 1521 1073
rect 1563 1065 1630 1073
rect 1673 1066 1740 1074
rect 1782 1065 1849 1073
rect 11 1004 46 1009
rect 938 998 1865 1021
rect 910 997 1865 998
rect 909 993 1865 997
rect 1785 986 1865 993
rect -34 878 30 893
rect -34 670 4 878
rect 1828 783 1865 986
rect 1790 770 1865 783
rect 1795 745 1807 753
rect 1790 727 1807 733
rect -34 654 30 670
rect -34 524 4 654
rect 1828 555 1865 770
rect 1790 547 1865 555
rect -34 513 30 524
rect -34 385 4 513
rect 1828 456 1865 547
rect 1787 443 1865 456
rect -34 369 30 385
rect -34 237 4 369
rect 1828 311 1865 443
rect 1790 295 1865 311
rect 1790 267 1798 277
rect -34 220 30 237
rect -34 36 4 220
rect 1790 123 1798 131
rect 1828 110 1865 295
rect 1790 94 1865 110
rect -34 20 31 36
rect 1828 19 1865 94
rect 88 -21 155 -13
rect 201 -19 268 -11
rect 309 -18 376 -10
rect 420 -18 487 -10
rect 532 -18 599 -10
rect 642 -17 709 -9
rect 754 -16 821 -8
rect 861 -15 928 -7
rect 969 -17 1036 -9
rect 1081 -16 1148 -8
rect 1192 -16 1259 -8
rect 1301 -15 1368 -7
rect 1411 -14 1478 -6
rect 1521 -14 1588 -6
rect 1631 -16 1698 -8
rect 1741 -17 1808 -9
<< metal2 >>
rect 43 1823 49 1856
rect 153 1823 159 1859
rect 263 1823 269 1856
rect 373 1823 379 1856
rect 483 1823 489 1856
rect 593 1823 599 1856
rect 703 1823 709 1856
rect 813 1823 819 1856
rect 925 1635 1936 1644
rect 1912 1625 1935 1635
rect 925 1617 997 1623
rect 1911 1504 1935 1625
rect 925 1446 1976 1453
rect 918 1316 1026 1324
rect 948 1198 956 1316
rect 1005 1072 1011 1073
rect 1115 1072 1121 1073
rect 1005 1064 1006 1072
rect 1115 1064 1117 1072
rect 1225 1071 1231 1073
rect 1005 994 1011 1064
rect 1115 994 1121 1064
rect 1225 1063 1227 1071
rect 1335 1066 1337 1073
rect 1225 994 1231 1063
rect 1335 994 1341 1066
rect 1445 1065 1448 1073
rect 1555 1065 1557 1073
rect 1665 1066 1667 1073
rect 1445 994 1451 1065
rect 1555 994 1561 1065
rect 1665 994 1671 1066
rect 1774 1065 1776 1073
rect 1774 994 1780 1065
rect 1812 745 1825 753
rect 1812 727 1823 733
rect 1790 493 1815 501
rect 1790 466 1814 469
rect 1794 462 1814 466
rect 1912 277 1935 1412
rect 1806 267 1937 277
rect 1954 133 1976 1446
rect 1803 131 1995 133
rect 1804 124 1995 131
rect 81 -13 94 20
rect 81 -21 82 -13
rect 88 -21 94 -13
rect 191 -11 204 20
rect 191 -19 195 -11
rect 201 -19 204 -11
rect 191 -21 204 -19
rect 301 -10 314 20
rect 301 -18 303 -10
rect 309 -18 314 -10
rect 301 -21 314 -18
rect 411 -10 424 20
rect 411 -18 414 -10
rect 420 -18 424 -10
rect 411 -21 424 -18
rect 521 -10 534 20
rect 521 -18 526 -10
rect 532 -18 534 -10
rect 521 -21 534 -18
rect 631 -9 644 20
rect 631 -17 636 -9
rect 642 -17 644 -9
rect 631 -21 644 -17
rect 741 -8 754 20
rect 741 -16 748 -8
rect 741 -21 754 -16
rect 851 -7 864 20
rect 851 -15 855 -7
rect 861 -15 864 -7
rect 851 -21 864 -15
rect 961 -9 974 20
rect 961 -17 963 -9
rect 969 -17 974 -9
rect 961 -21 974 -17
rect 1071 -8 1084 20
rect 1071 -16 1075 -8
rect 1081 -16 1084 -8
rect 1071 -21 1084 -16
rect 1181 -8 1194 20
rect 1181 -16 1186 -8
rect 1192 -16 1194 -8
rect 1181 -21 1194 -16
rect 1291 -7 1304 20
rect 1291 -15 1295 -7
rect 1301 -15 1304 -7
rect 1291 -21 1304 -15
rect 1401 -6 1414 20
rect 1401 -14 1405 -6
rect 1411 -14 1414 -6
rect 1401 -21 1414 -14
rect 1511 -6 1524 20
rect 1511 -14 1515 -6
rect 1521 -14 1524 -6
rect 1511 -21 1524 -14
rect 1621 -8 1634 20
rect 1621 -16 1625 -8
rect 1631 -16 1634 -8
rect 1621 -21 1634 -16
rect 1731 -9 1744 20
rect 1731 -17 1735 -9
rect 1741 -17 1744 -9
rect 1731 -21 1744 -17
<< ntransistor >>
rect 918 1199 928 1201
<< ptransistor >>
rect 917 1155 935 1157
<< polycontact >>
rect 910 1635 915 1643
rect 942 1178 948 1184
rect 1790 745 1795 753
<< ndcontact >>
rect 918 1203 928 1209
rect 918 1191 928 1197
<< pdcontact >>
rect 917 1159 935 1166
rect 917 1146 935 1153
<< m2contact >>
rect 43 1856 49 1864
rect 153 1859 159 1867
rect 263 1856 269 1864
rect 373 1856 379 1864
rect 483 1856 489 1864
rect 593 1856 599 1864
rect 703 1856 709 1864
rect 813 1856 819 1864
rect 920 1635 925 1643
rect 920 1617 925 1623
rect 919 1446 925 1454
rect 1911 1484 1937 1504
rect 910 1316 918 1324
rect 1912 1412 1935 1424
rect 948 1190 956 1198
rect 1006 1064 1012 1072
rect 1117 1064 1123 1072
rect 1227 1063 1233 1071
rect 1337 1066 1343 1074
rect 1448 1065 1454 1073
rect 1557 1065 1563 1073
rect 1667 1066 1673 1074
rect 1776 1065 1782 1073
rect 46 1004 50 1009
rect 1807 745 1812 753
rect 1807 727 1812 733
rect 1790 462 1794 466
rect 1798 267 1806 277
rect 1798 123 1804 131
rect 82 -21 88 -13
rect 195 -19 201 -11
rect 303 -18 309 -10
rect 414 -18 420 -10
rect 526 -18 532 -10
rect 636 -17 642 -9
rect 748 -16 754 -8
rect 855 -15 861 -7
rect 963 -17 969 -9
rect 1075 -16 1081 -8
rect 1186 -16 1192 -8
rect 1295 -15 1301 -7
rect 1405 -14 1411 -6
rect 1515 -14 1521 -6
rect 1625 -16 1631 -8
rect 1735 -17 1741 -9
use datapathL  datapathL_0 ../cells
array 0 7 110 0 0 1803
timestamp 1428628260
transform 1 0 30 0 1 562
box 0 -542 110 1261
use datapathS  datapathS_0 ../cells
array 0 7 110 0 0 974
timestamp 1428625343
transform 1 0 910 0 1 562
box 0 -542 110 432
<< labels >>
rlabel metal2 1790 495 1815 499 0 INBIT
rlabel metal1 -34 20 4 1822 0 Vdd
rlabel metal1 1828 19 1865 1021 0 GND
rlabel metal2 925 1617 997 1623 0 CLKLD
rlabel metal2 925 1635 1936 1644 0 CLK
rlabel metal2 918 1316 1026 1324 0 ADDSUB
rlabel space 1774 988 1780 1073 1 DIVIDEND_0
rlabel space 1665 988 1671 1073 1 DIVIDEND_1
rlabel space 1555 988 1561 1073 1 DIVIDEND_2
rlabel space 1445 988 1451 1073 1 DIVIDEND_3
rlabel space 1335 988 1341 1073 1 DIVIDEND_4
rlabel space 1225 988 1231 1073 1 DIVIDEND_5
rlabel space 1115 988 1121 1073 1 DIVIDEND_6
rlabel space 1005 988 1011 1073 1 DIVIDEND_7
rlabel metal2 1794 462 1814 469 0 SHIFT
rlabel metal2 1812 727 1823 733 0 S1
rlabel metal2 1812 745 1825 753 0 S0
rlabel metal1 11 1004 46 1009 0 SIGN
rlabel metal1 819 1856 886 1864 1 DIVISOR_0
rlabel metal1 709 1856 776 1864 1 DIVISOR_1
rlabel metal1 599 1856 666 1864 1 DIVISOR_2
rlabel metal1 489 1856 556 1864 1 DIVISOR_3
rlabel metal1 379 1856 446 1864 1 DIVISOR_4
rlabel metal1 269 1856 336 1864 1 DIVISOR_5
rlabel metal1 159 1859 226 1867 5 DIVISOR_6
rlabel metal1 49 1856 116 1864 1 DIVISOR_7
rlabel metal1 1782 1065 1849 1073 1 DIVIDEND_0
rlabel metal1 1673 1066 1740 1074 1 DIVIDEND_1
rlabel metal1 1563 1065 1630 1073 1 DIVIDEND_2
rlabel metal1 1454 1065 1521 1073 1 DIVIDEND_3
rlabel metal1 1343 1066 1410 1074 1 DIVIDEND_4
rlabel metal1 1233 1063 1300 1071 1 DIVIDEND_5
rlabel metal1 1123 1064 1190 1072 1 DIVIDEND_6
rlabel metal1 1012 1064 1079 1072 1 DIVIDEND_7
rlabel metal1 1741 -17 1808 -9 1 REM_0
rlabel metal1 1631 -16 1698 -8 1 REM_1
rlabel metal1 1521 -14 1588 -6 1 REM_2
rlabel metal1 1411 -14 1478 -6 1 REM_3
rlabel metal1 1301 -15 1368 -7 1 REM_4
rlabel metal1 1192 -16 1259 -8 1 REM_5
rlabel metal1 1081 -16 1148 -8 1 REM_6
rlabel metal1 969 -17 1036 -9 1 REM_7
rlabel metal1 861 -15 928 -7 1 REM_8
rlabel metal1 754 -16 821 -8 1 REM_9
rlabel metal1 642 -17 709 -9 1 REM_10
rlabel metal1 532 -18 599 -10 1 REM_11
rlabel metal1 420 -18 487 -10 1 REM_12
rlabel metal1 309 -18 376 -10 1 REM_13
rlabel metal1 201 -19 268 -11 1 REM_14
rlabel metal1 88 -21 155 -13 1 REM_15
rlabel metal2 1954 124 1976 1453 0 RST
<< end >>
