magic
tech scmos
timestamp 1428807341
<< pwell >>
rect 125 322 139 356
rect 123 177 139 233
rect 452 111 475 140
rect 385 71 475 111
rect 123 -24 139 58
rect 385 -44 475 -4
rect 452 -73 475 -44
rect 226 -143 388 -115
<< nwell >>
rect 123 239 139 316
rect 123 64 139 171
rect 385 115 449 145
rect 385 0 475 67
rect 123 -78 139 -30
rect 385 -65 448 -48
rect 378 -70 448 -65
rect 226 -78 448 -70
rect 226 -80 397 -78
rect 226 -111 388 -80
<< polysilicon >>
rect 449 139 462 141
rect 449 138 451 139
rect 460 138 462 139
rect 406 134 408 138
rect 416 134 418 138
rect 426 134 428 138
rect 436 134 438 138
rect 406 116 408 118
rect 397 111 408 116
rect 416 115 418 118
rect 417 111 418 115
rect 406 108 408 111
rect 416 108 418 111
rect 426 108 428 118
rect 436 108 438 118
rect 406 96 408 98
rect 416 96 418 98
rect 406 84 408 86
rect 416 84 418 86
rect 426 84 428 98
rect 436 84 438 98
rect 460 96 462 98
rect 445 86 456 88
rect 406 64 408 74
rect 416 72 418 74
rect 426 72 428 74
rect 416 70 428 72
rect 416 64 418 70
rect 426 64 428 70
rect 436 64 438 74
rect 445 67 447 86
rect 454 84 456 86
rect 464 84 466 86
rect 454 64 456 74
rect 464 64 466 74
rect 406 38 408 44
rect 416 42 418 44
rect 398 36 408 38
rect 398 30 400 36
rect 426 30 428 44
rect 398 26 399 30
rect 427 26 428 30
rect 398 23 400 26
rect 416 23 418 25
rect 426 23 428 26
rect 436 30 438 44
rect 454 42 456 44
rect 464 30 466 44
rect 436 26 437 30
rect 465 26 466 30
rect 436 23 438 26
rect 446 23 448 25
rect 464 23 466 26
rect 398 -7 400 3
rect 416 0 418 3
rect 407 -4 418 0
rect 416 -7 418 -4
rect 426 -7 428 3
rect 436 -7 438 3
rect 446 0 448 3
rect 446 -4 457 0
rect 446 -7 448 -4
rect 464 -7 466 3
rect 398 -19 400 -17
rect 416 -19 418 -17
rect 416 -31 418 -29
rect 426 -31 428 -17
rect 436 -31 438 -17
rect 446 -19 448 -17
rect 464 -19 466 -17
rect 460 -31 462 -29
rect 416 -44 418 -41
rect 417 -48 418 -44
rect 416 -52 418 -48
rect 426 -52 428 -41
rect 436 -52 438 -41
rect 416 -78 418 -68
rect 199 -80 244 -78
rect 199 -81 202 -80
rect 242 -81 244 -80
rect 252 -81 254 -79
rect 262 -81 264 -79
rect 272 -81 274 -79
rect 309 -80 347 -78
rect 309 -81 312 -80
rect 345 -81 347 -80
rect 355 -81 357 -79
rect 365 -81 367 -79
rect 375 -81 377 -79
rect 426 -81 428 -68
rect 436 -88 438 -68
rect 449 -72 451 -71
rect 460 -72 462 -71
rect 449 -74 462 -72
rect 429 -91 438 -88
rect 242 -118 244 -108
rect 252 -111 254 -108
rect 253 -115 254 -111
rect 252 -118 254 -115
rect 262 -118 264 -108
rect 272 -118 274 -108
rect 345 -118 347 -108
rect 355 -111 357 -108
rect 356 -115 357 -111
rect 355 -118 357 -115
rect 365 -118 367 -108
rect 375 -118 377 -108
rect 242 -135 244 -133
rect 252 -134 254 -133
rect 262 -134 264 -133
rect 272 -134 274 -133
rect 252 -136 274 -134
rect 345 -135 347 -133
rect 355 -134 357 -133
rect 365 -134 367 -133
rect 375 -134 377 -133
rect 355 -136 377 -134
<< ndiffusion >>
rect 404 98 406 108
rect 408 98 410 108
rect 414 98 416 108
rect 418 98 426 108
rect 428 98 436 108
rect 438 98 440 108
rect 458 98 460 138
rect 462 98 464 138
rect 404 74 406 84
rect 408 74 416 84
rect 418 74 420 84
rect 424 74 426 84
rect 428 74 430 84
rect 434 74 436 84
rect 438 74 440 84
rect 452 74 454 84
rect 456 74 458 84
rect 462 74 464 84
rect 466 74 468 84
rect 396 -17 398 -7
rect 400 -17 402 -7
rect 414 -17 416 -7
rect 418 -17 420 -7
rect 424 -17 426 -7
rect 428 -17 430 -7
rect 434 -17 436 -7
rect 438 -17 440 -7
rect 444 -17 446 -7
rect 448 -17 450 -7
rect 462 -17 464 -7
rect 466 -17 468 -7
rect 414 -41 416 -31
rect 418 -41 426 -31
rect 428 -41 436 -31
rect 438 -41 440 -31
rect 458 -71 460 -31
rect 462 -71 464 -31
rect 240 -133 242 -118
rect 244 -133 246 -118
rect 250 -133 252 -118
rect 254 -133 256 -118
rect 260 -133 262 -118
rect 264 -133 266 -118
rect 270 -133 272 -118
rect 274 -133 276 -118
rect 343 -133 345 -118
rect 347 -133 349 -118
rect 353 -133 355 -118
rect 357 -133 359 -118
rect 363 -133 365 -118
rect 367 -133 369 -118
rect 373 -133 375 -118
rect 377 -133 379 -118
<< pdiffusion >>
rect 404 118 406 134
rect 408 118 410 134
rect 414 118 416 134
rect 418 118 420 134
rect 424 118 426 134
rect 428 118 430 134
rect 434 118 436 134
rect 438 118 440 134
rect 404 44 406 64
rect 408 44 410 64
rect 414 44 416 64
rect 418 44 420 64
rect 424 44 426 64
rect 428 44 436 64
rect 438 44 440 64
rect 452 44 454 64
rect 456 44 458 64
rect 462 44 464 64
rect 466 44 468 64
rect 396 3 398 23
rect 400 3 402 23
rect 414 3 416 23
rect 418 3 420 23
rect 424 3 426 23
rect 428 3 430 23
rect 434 3 436 23
rect 438 3 440 23
rect 444 3 446 23
rect 448 3 450 23
rect 462 3 464 23
rect 466 3 468 23
rect 414 -68 416 -52
rect 418 -68 420 -52
rect 424 -68 426 -52
rect 428 -68 430 -52
rect 434 -68 436 -52
rect 438 -68 440 -52
rect 240 -108 242 -81
rect 244 -108 246 -81
rect 250 -108 252 -81
rect 254 -108 256 -81
rect 260 -108 262 -81
rect 264 -108 266 -81
rect 270 -108 272 -81
rect 274 -108 276 -81
rect 343 -108 345 -81
rect 347 -108 349 -81
rect 353 -108 355 -81
rect 357 -108 359 -81
rect 363 -108 365 -81
rect 367 -108 369 -81
rect 373 -108 375 -81
rect 377 -108 379 -81
<< metal1 >>
rect 128 345 135 362
rect 128 271 134 287
rect 128 197 134 213
rect 347 169 376 179
rect 368 163 376 169
rect 358 157 365 161
rect 354 145 358 149
rect 361 152 365 157
rect 368 155 532 163
rect 361 148 424 152
rect 354 142 360 145
rect 128 123 134 139
rect 356 138 360 142
rect 369 141 386 145
rect 396 141 413 145
rect 356 134 369 138
rect 410 134 414 141
rect 360 122 369 134
rect 360 118 393 122
rect 420 134 424 148
rect 434 141 475 145
rect 430 134 434 141
rect 447 133 451 134
rect 444 118 454 123
rect 400 115 404 118
rect 420 115 424 118
rect 440 115 454 118
rect 393 110 397 111
rect 349 102 373 110
rect 400 111 413 115
rect 420 111 454 115
rect 400 108 404 111
rect 440 108 454 111
rect 349 33 357 102
rect 444 98 454 108
rect 471 125 475 129
rect 471 102 475 106
rect 410 95 414 98
rect 464 95 468 98
rect 381 94 475 95
rect 381 88 397 94
rect 420 88 457 94
rect 471 88 475 94
rect 381 87 475 88
rect 420 84 424 87
rect 440 84 444 87
rect 458 84 462 87
rect 400 71 404 74
rect 430 71 434 74
rect 448 71 452 74
rect 400 67 410 71
rect 434 67 441 71
rect 410 64 414 67
rect 440 64 444 67
rect 448 64 452 67
rect 468 71 472 74
rect 468 67 475 71
rect 468 64 472 67
rect 400 41 404 44
rect 420 41 424 44
rect 458 41 462 44
rect 369 40 475 41
rect 369 33 442 40
rect 463 33 475 40
rect 129 25 134 33
rect 348 25 357 33
rect 392 23 396 33
rect 403 26 409 30
rect 422 26 423 30
rect 430 23 434 33
rect 441 26 442 30
rect 460 26 461 30
rect 468 23 472 33
rect 128 -4 134 12
rect 348 -4 373 12
rect 406 3 407 23
rect 403 0 407 3
rect 410 0 414 3
rect 450 0 454 3
rect 410 -4 420 0
rect 403 -7 407 -4
rect 420 -7 424 -4
rect 444 -4 454 0
rect 457 3 458 23
rect 457 0 461 3
rect 472 -4 475 0
rect 440 -7 444 -4
rect 457 -7 461 -4
rect 406 -17 407 -7
rect 457 -17 458 -7
rect 392 -20 396 -17
rect 410 -20 414 -17
rect 430 -20 434 -17
rect 450 -20 454 -17
rect 468 -20 472 -17
rect 381 -21 475 -20
rect 381 -27 395 -21
rect 420 -27 475 -21
rect 381 -28 475 -27
rect 410 -31 414 -28
rect 464 -31 468 -28
rect 444 -41 454 -31
rect 440 -44 454 -41
rect 397 -48 413 -44
rect 424 -48 454 -44
rect 420 -52 424 -48
rect 440 -51 454 -48
rect 440 -52 444 -51
rect 128 -78 134 -62
rect 346 -78 361 -62
rect 447 -67 451 -66
rect 410 -74 414 -68
rect 430 -74 434 -68
rect 471 -39 475 -35
rect 369 -78 387 -74
rect 406 -78 475 -74
rect 246 -81 250 -78
rect 266 -81 270 -78
rect 349 -81 353 -78
rect 369 -81 373 -78
rect 197 -85 198 -81
rect 215 -136 223 -86
rect 307 -85 308 -81
rect 280 -94 281 -90
rect 236 -111 240 -108
rect 256 -111 260 -108
rect 276 -111 280 -108
rect 236 -115 249 -111
rect 256 -115 280 -111
rect 236 -118 240 -115
rect 256 -118 260 -115
rect 276 -118 280 -115
rect 383 -85 425 -81
rect 423 -90 425 -88
rect 424 -92 425 -90
rect 424 -94 427 -92
rect 339 -111 343 -108
rect 359 -111 363 -108
rect 379 -111 383 -108
rect 339 -115 352 -111
rect 359 -115 383 -111
rect 524 -115 532 155
rect 339 -118 343 -115
rect 359 -118 363 -115
rect 379 -118 383 -115
rect 246 -136 250 -133
rect 266 -136 270 -133
rect 349 -136 353 -133
rect 369 -136 373 -133
rect 215 -141 297 -136
rect 321 -141 393 -136
<< metal2 >>
rect 148 363 366 366
rect 148 358 154 363
rect 258 352 358 358
rect 354 161 358 352
rect 362 153 366 363
rect 358 149 366 153
rect 373 151 540 159
rect 363 130 369 141
rect 361 41 369 130
rect 373 110 381 151
rect 417 141 430 145
rect 385 129 447 130
rect 385 126 451 129
rect 184 -81 197 -77
rect 233 -81 241 -1
rect 361 -62 369 33
rect 373 12 381 87
rect 373 -20 381 -4
rect 385 -52 389 126
rect 464 122 471 125
rect 397 118 405 122
rect 393 -44 397 106
rect 401 -39 405 118
rect 410 121 471 122
rect 410 118 468 121
rect 410 71 414 118
rect 430 98 471 102
rect 430 71 434 98
rect 448 63 475 67
rect 409 34 446 38
rect 409 30 413 34
rect 442 30 446 34
rect 418 22 422 26
rect 456 22 460 26
rect 418 18 460 22
rect 444 -4 468 0
rect 420 -31 424 -4
rect 420 -35 471 -31
rect 401 -43 424 -39
rect 420 -44 424 -43
rect 385 -56 451 -52
rect 223 -86 241 -81
rect 294 -81 307 -76
rect 447 -62 451 -56
rect 285 -94 420 -90
<< ntransistor >>
rect 406 98 408 108
rect 416 98 418 108
rect 426 98 428 108
rect 436 98 438 108
rect 460 98 462 138
rect 406 74 408 84
rect 416 74 418 84
rect 426 74 428 84
rect 436 74 438 84
rect 454 74 456 84
rect 464 74 466 84
rect 398 -17 400 -7
rect 416 -17 418 -7
rect 426 -17 428 -7
rect 436 -17 438 -7
rect 446 -17 448 -7
rect 464 -17 466 -7
rect 416 -41 418 -31
rect 426 -41 428 -31
rect 436 -41 438 -31
rect 460 -71 462 -31
rect 242 -133 244 -118
rect 252 -133 254 -118
rect 262 -133 264 -118
rect 272 -133 274 -118
rect 345 -133 347 -118
rect 355 -133 357 -118
rect 365 -133 367 -118
rect 375 -133 377 -118
<< ptransistor >>
rect 406 118 408 134
rect 416 118 418 134
rect 426 118 428 134
rect 436 118 438 134
rect 406 44 408 64
rect 416 44 418 64
rect 426 44 428 64
rect 436 44 438 64
rect 454 44 456 64
rect 464 44 466 64
rect 398 3 400 23
rect 416 3 418 23
rect 426 3 428 23
rect 436 3 438 23
rect 446 3 448 23
rect 464 3 466 23
rect 416 -68 418 -52
rect 426 -68 428 -52
rect 436 -68 438 -52
rect 242 -108 244 -81
rect 252 -108 254 -81
rect 262 -108 264 -81
rect 272 -108 274 -81
rect 345 -108 347 -81
rect 355 -108 357 -81
rect 365 -108 367 -81
rect 375 -108 377 -81
<< polycontact >>
rect 447 134 451 138
rect 393 111 397 115
rect 413 111 417 115
rect 441 67 445 71
rect 399 26 403 30
rect 423 26 427 30
rect 437 26 441 30
rect 461 26 465 30
rect 403 -4 407 0
rect 457 -4 461 0
rect 413 -48 417 -44
rect 198 -85 202 -81
rect 308 -85 312 -81
rect 425 -85 429 -81
rect 447 -71 451 -67
rect 425 -92 429 -88
rect 249 -115 253 -111
rect 352 -115 356 -111
<< ndcontact >>
rect 400 98 404 108
rect 410 98 414 108
rect 440 98 444 108
rect 454 98 458 138
rect 464 98 468 138
rect 400 74 404 84
rect 420 74 424 84
rect 430 74 434 84
rect 440 74 444 84
rect 448 74 452 84
rect 458 74 462 84
rect 468 74 472 84
rect 392 -17 396 -7
rect 402 -17 406 -7
rect 410 -17 414 -7
rect 420 -17 424 -7
rect 430 -17 434 -7
rect 440 -17 444 -7
rect 450 -17 454 -7
rect 458 -17 462 -7
rect 468 -17 472 -7
rect 410 -41 414 -31
rect 440 -41 444 -31
rect 454 -71 458 -31
rect 464 -71 468 -31
rect 236 -133 240 -118
rect 246 -133 250 -118
rect 256 -133 260 -118
rect 266 -133 270 -118
rect 276 -133 280 -118
rect 339 -133 343 -118
rect 349 -133 353 -118
rect 359 -133 363 -118
rect 369 -133 373 -118
rect 379 -133 383 -118
<< pdcontact >>
rect 400 118 404 134
rect 410 118 414 134
rect 420 118 424 134
rect 430 118 434 134
rect 440 118 444 134
rect 400 44 404 64
rect 410 44 414 64
rect 420 44 424 64
rect 440 44 444 64
rect 448 44 452 64
rect 458 44 462 64
rect 468 44 472 64
rect 392 3 396 23
rect 402 3 406 23
rect 410 3 414 23
rect 420 3 424 23
rect 430 3 434 23
rect 440 3 444 23
rect 450 3 454 23
rect 458 3 462 23
rect 468 3 472 23
rect 410 -68 414 -52
rect 420 -68 424 -52
rect 430 -68 434 -52
rect 440 -68 444 -52
rect 236 -108 240 -81
rect 246 -108 250 -81
rect 256 -108 260 -81
rect 266 -108 270 -81
rect 276 -108 280 -81
rect 339 -108 343 -81
rect 349 -108 353 -81
rect 359 -108 363 -81
rect 369 -108 373 -81
rect 379 -108 383 -81
<< m2contact >>
rect 354 157 358 161
rect 354 149 358 153
rect 363 141 369 145
rect 413 141 417 145
rect 393 118 397 122
rect 430 141 434 145
rect 447 129 451 133
rect 373 102 381 110
rect 393 106 397 110
rect 471 121 475 125
rect 471 98 475 102
rect 373 87 381 95
rect 410 67 414 71
rect 430 67 434 71
rect 448 67 452 71
rect 361 33 369 41
rect 409 26 413 30
rect 418 26 422 30
rect 442 26 446 30
rect 456 26 460 30
rect 233 -1 241 8
rect 373 -4 381 12
rect 420 -4 424 0
rect 440 -4 444 0
rect 468 -4 472 0
rect 373 -28 381 -20
rect 393 -48 397 -44
rect 420 -48 424 -44
rect 361 -78 369 -62
rect 447 -66 451 -62
rect 471 -35 475 -31
rect 184 -85 197 -81
rect 215 -86 223 -81
rect 294 -85 307 -81
rect 281 -94 285 -90
rect 420 -94 424 -90
rect 540 151 548 159
<< psubstratepcontact >>
rect 397 88 420 94
rect 457 88 471 94
rect 395 -27 420 -21
rect 297 -141 321 -136
<< nsubstratencontact >>
rect 386 138 396 145
rect 442 33 463 40
rect 387 -78 406 -74
use rego  rego_0 ../cells
timestamp 1428793378
transform 1 0 133 0 1 82
box 0 -160 110 279
use rego  rego_1
timestamp 1428793378
transform 1 0 243 0 1 82
box 0 -160 110 279
<< labels >>
rlabel space 361 41 369 141 3 Vdd
rlabel metal2 385 -56 451 -52 1 start
rlabel metal1 420 -48 444 -44 1 nextSB1
rlabel metal1 471 -39 475 -35 1 inbit
rlabel metal1 471 125 475 129 1 shift
rlabel metal1 471 102 475 106 1 load
rlabel metal1 420 111 444 115 1 nextSB0
rlabel metal2 374 -28 380 95 3 Gnd
rlabel polysilicon 436 -81 438 -71 1 SB1
rlabel polysilicon 426 -81 428 -71 1 SB0
rlabel metal1 397 -48 413 -44 1 sign
rlabel metal1 472 -4 475 0 7 add
rlabel metal2 448 63 475 67 1 sel0
rlabel metal1 468 64 472 74 1 sel1
rlabel metal1 420 136 424 152 1 nextSB0
rlabel metal2 401 -43 424 -39 1 nextSB1
rlabel metal1 524 -115 532 163 1 clk
<< end >>
