magic
tech scmos
timestamp 1428890255
<< pwell >>
rect 993 1566 1103 1570
rect 993 1561 1229 1566
rect 993 1548 1653 1561
rect 993 1545 1229 1548
rect 993 1542 1101 1545
rect 1425 1370 1438 1380
rect 1747 1362 1770 1383
rect 902 1185 926 1267
rect 1421 1166 1446 1184
rect 1727 986 1773 1068
rect 1882 23 1897 2023
rect 1939 23 1965 2023
<< nwell >>
rect 1748 1387 1770 1418
rect 903 1121 926 1181
rect 909 1116 926 1121
rect 1711 1071 1773 1117
rect 1901 23 1935 2023
rect 1969 23 1988 2023
<< polysilicon >>
rect 1874 2022 1901 2024
rect 1897 2015 1901 2022
rect 1935 2023 1969 2024
rect 1939 2022 1969 2023
rect 1888 2013 1890 2015
rect 1894 2013 1904 2015
rect 1912 2013 1914 2015
rect 1888 2005 1890 2007
rect 1894 2006 1897 2007
rect 1901 2006 1904 2007
rect 1894 2005 1904 2006
rect 1912 2005 1914 2007
rect 1922 2014 1924 2016
rect 1932 2015 1942 2016
rect 1932 2014 1935 2015
rect 1939 2014 1942 2015
rect 1946 2014 1948 2016
rect 1965 2015 1969 2022
rect 1922 2006 1924 2008
rect 1932 2006 1942 2008
rect 1946 2006 1948 2008
rect 1956 2013 1958 2015
rect 1962 2013 1972 2015
rect 1980 2013 1982 2015
rect 1897 1990 1901 1998
rect 1935 1998 1939 2006
rect 1956 2005 1958 2007
rect 1962 2006 1965 2007
rect 1969 2006 1972 2007
rect 1962 2005 1972 2006
rect 1980 2005 1982 2007
rect 1888 1988 1890 1990
rect 1894 1988 1904 1990
rect 1912 1988 1914 1990
rect 1888 1980 1890 1982
rect 1894 1981 1897 1982
rect 1901 1981 1904 1982
rect 1894 1980 1904 1981
rect 1912 1980 1914 1982
rect 1922 1989 1924 1991
rect 1932 1990 1942 1991
rect 1932 1989 1935 1990
rect 1939 1989 1942 1990
rect 1946 1989 1948 1991
rect 1965 1990 1969 1998
rect 1922 1981 1924 1983
rect 1932 1981 1942 1983
rect 1946 1981 1948 1983
rect 1956 1988 1958 1990
rect 1962 1988 1972 1990
rect 1980 1988 1982 1990
rect 1897 1965 1901 1973
rect 1935 1973 1939 1981
rect 1956 1980 1958 1982
rect 1962 1981 1965 1982
rect 1969 1981 1972 1982
rect 1962 1980 1972 1981
rect 1980 1980 1982 1982
rect 1888 1963 1890 1965
rect 1894 1963 1904 1965
rect 1912 1963 1914 1965
rect 1888 1955 1890 1957
rect 1894 1956 1897 1957
rect 1901 1956 1904 1957
rect 1894 1955 1904 1956
rect 1912 1955 1914 1957
rect 1922 1964 1924 1966
rect 1932 1965 1942 1966
rect 1932 1964 1935 1965
rect 1939 1964 1942 1965
rect 1946 1964 1948 1966
rect 1965 1965 1969 1973
rect 1922 1956 1924 1958
rect 1932 1956 1942 1958
rect 1946 1956 1948 1958
rect 1956 1963 1958 1965
rect 1962 1963 1972 1965
rect 1980 1963 1982 1965
rect 1897 1940 1901 1948
rect 1935 1948 1939 1956
rect 1956 1955 1958 1957
rect 1962 1956 1965 1957
rect 1969 1956 1972 1957
rect 1962 1955 1972 1956
rect 1980 1955 1982 1957
rect 1888 1938 1890 1940
rect 1894 1938 1904 1940
rect 1912 1938 1914 1940
rect 1888 1930 1890 1932
rect 1894 1931 1897 1932
rect 1901 1931 1904 1932
rect 1894 1930 1904 1931
rect 1912 1930 1914 1932
rect 1922 1939 1924 1941
rect 1932 1940 1942 1941
rect 1932 1939 1935 1940
rect 1939 1939 1942 1940
rect 1946 1939 1948 1941
rect 1965 1940 1969 1948
rect 1922 1931 1924 1933
rect 1932 1931 1942 1933
rect 1946 1931 1948 1933
rect 1956 1938 1958 1940
rect 1962 1938 1972 1940
rect 1980 1938 1982 1940
rect 1897 1915 1901 1923
rect 1935 1923 1939 1931
rect 1956 1930 1958 1932
rect 1962 1931 1965 1932
rect 1969 1931 1972 1932
rect 1962 1930 1972 1931
rect 1980 1930 1982 1932
rect 1888 1913 1890 1915
rect 1894 1913 1904 1915
rect 1912 1913 1914 1915
rect 1888 1905 1890 1907
rect 1894 1906 1897 1907
rect 1901 1906 1904 1907
rect 1894 1905 1904 1906
rect 1912 1905 1914 1907
rect 1922 1914 1924 1916
rect 1932 1915 1942 1916
rect 1932 1914 1935 1915
rect 1939 1914 1942 1915
rect 1946 1914 1948 1916
rect 1965 1915 1969 1923
rect 1922 1906 1924 1908
rect 1932 1906 1942 1908
rect 1946 1906 1948 1908
rect 1956 1913 1958 1915
rect 1962 1913 1972 1915
rect 1980 1913 1982 1915
rect 1897 1890 1901 1898
rect 1935 1898 1939 1906
rect 1956 1905 1958 1907
rect 1962 1906 1965 1907
rect 1969 1906 1972 1907
rect 1962 1905 1972 1906
rect 1980 1905 1982 1907
rect 1888 1888 1890 1890
rect 1894 1888 1904 1890
rect 1912 1888 1914 1890
rect 1888 1880 1890 1882
rect 1894 1881 1897 1882
rect 1901 1881 1904 1882
rect 1894 1880 1904 1881
rect 1912 1880 1914 1882
rect 1922 1889 1924 1891
rect 1932 1890 1942 1891
rect 1932 1889 1935 1890
rect 1939 1889 1942 1890
rect 1946 1889 1948 1891
rect 1965 1890 1969 1898
rect 1922 1881 1924 1883
rect 1932 1881 1942 1883
rect 1946 1881 1948 1883
rect 1956 1888 1958 1890
rect 1962 1888 1972 1890
rect 1980 1888 1982 1890
rect 1897 1865 1901 1873
rect 1935 1873 1939 1881
rect 1956 1880 1958 1882
rect 1962 1881 1965 1882
rect 1969 1881 1972 1882
rect 1962 1880 1972 1881
rect 1980 1880 1982 1882
rect 1888 1863 1890 1865
rect 1894 1863 1904 1865
rect 1912 1863 1914 1865
rect 1888 1855 1890 1857
rect 1894 1856 1897 1857
rect 1901 1856 1904 1857
rect 1894 1855 1904 1856
rect 1912 1855 1914 1857
rect 1922 1864 1924 1866
rect 1932 1865 1942 1866
rect 1932 1864 1935 1865
rect 1939 1864 1942 1865
rect 1946 1864 1948 1866
rect 1965 1865 1969 1873
rect 1922 1856 1924 1858
rect 1932 1856 1942 1858
rect 1946 1856 1948 1858
rect 1956 1863 1958 1865
rect 1962 1863 1972 1865
rect 1980 1863 1982 1865
rect 1897 1840 1901 1848
rect 1935 1848 1939 1856
rect 1956 1855 1958 1857
rect 1962 1856 1965 1857
rect 1969 1856 1972 1857
rect 1962 1855 1972 1856
rect 1980 1855 1982 1857
rect 1888 1838 1890 1840
rect 1894 1838 1904 1840
rect 1912 1838 1914 1840
rect 1888 1830 1890 1832
rect 1894 1831 1897 1832
rect 1901 1831 1904 1832
rect 1894 1830 1904 1831
rect 1912 1830 1914 1832
rect 1922 1839 1924 1841
rect 1932 1840 1942 1841
rect 1932 1839 1935 1840
rect 1939 1839 1942 1840
rect 1946 1839 1948 1841
rect 1965 1840 1969 1848
rect 1922 1831 1924 1833
rect 1932 1831 1942 1833
rect 1946 1831 1948 1833
rect 1956 1838 1958 1840
rect 1962 1838 1972 1840
rect 1980 1838 1982 1840
rect 1897 1815 1901 1823
rect 1935 1823 1939 1831
rect 1956 1830 1958 1832
rect 1962 1831 1965 1832
rect 1969 1831 1972 1832
rect 1962 1830 1972 1831
rect 1980 1830 1982 1832
rect 1888 1813 1890 1815
rect 1894 1813 1904 1815
rect 1912 1813 1914 1815
rect 1888 1805 1890 1807
rect 1894 1806 1897 1807
rect 1901 1806 1904 1807
rect 1894 1805 1904 1806
rect 1912 1805 1914 1807
rect 1922 1814 1924 1816
rect 1932 1815 1942 1816
rect 1932 1814 1935 1815
rect 1939 1814 1942 1815
rect 1946 1814 1948 1816
rect 1965 1815 1969 1823
rect 1922 1806 1924 1808
rect 1932 1806 1942 1808
rect 1946 1806 1948 1808
rect 1956 1813 1958 1815
rect 1962 1813 1972 1815
rect 1980 1813 1982 1815
rect 1897 1790 1901 1798
rect 1935 1798 1939 1806
rect 1956 1805 1958 1807
rect 1962 1806 1965 1807
rect 1969 1806 1972 1807
rect 1962 1805 1972 1806
rect 1980 1805 1982 1807
rect 1888 1788 1890 1790
rect 1894 1788 1904 1790
rect 1912 1788 1914 1790
rect 1888 1780 1890 1782
rect 1894 1781 1897 1782
rect 1901 1781 1904 1782
rect 1894 1780 1904 1781
rect 1912 1780 1914 1782
rect 1922 1789 1924 1791
rect 1932 1790 1942 1791
rect 1932 1789 1935 1790
rect 1939 1789 1942 1790
rect 1946 1789 1948 1791
rect 1965 1790 1969 1798
rect 1922 1781 1924 1783
rect 1932 1781 1942 1783
rect 1946 1781 1948 1783
rect 1956 1788 1958 1790
rect 1962 1788 1972 1790
rect 1980 1788 1982 1790
rect 1897 1765 1901 1773
rect 1935 1773 1939 1781
rect 1956 1780 1958 1782
rect 1962 1781 1965 1782
rect 1969 1781 1972 1782
rect 1962 1780 1972 1781
rect 1980 1780 1982 1782
rect 1888 1763 1890 1765
rect 1894 1763 1904 1765
rect 1912 1763 1914 1765
rect 1888 1755 1890 1757
rect 1894 1756 1897 1757
rect 1901 1756 1904 1757
rect 1894 1755 1904 1756
rect 1912 1755 1914 1757
rect 1922 1764 1924 1766
rect 1932 1765 1942 1766
rect 1932 1764 1935 1765
rect 1939 1764 1942 1765
rect 1946 1764 1948 1766
rect 1965 1765 1969 1773
rect 1922 1756 1924 1758
rect 1932 1756 1942 1758
rect 1946 1756 1948 1758
rect 1956 1763 1958 1765
rect 1962 1763 1972 1765
rect 1980 1763 1982 1765
rect 1424 1670 1428 1744
rect 1897 1740 1901 1748
rect 1935 1748 1939 1756
rect 1956 1755 1958 1757
rect 1962 1756 1965 1757
rect 1969 1756 1972 1757
rect 1962 1755 1972 1756
rect 1980 1755 1982 1757
rect 1888 1738 1890 1740
rect 1894 1738 1904 1740
rect 1912 1738 1914 1740
rect 1888 1730 1890 1732
rect 1894 1731 1897 1732
rect 1901 1731 1904 1732
rect 1894 1730 1904 1731
rect 1912 1730 1914 1732
rect 1922 1739 1924 1741
rect 1932 1740 1942 1741
rect 1932 1739 1935 1740
rect 1939 1739 1942 1740
rect 1946 1739 1948 1741
rect 1965 1740 1969 1748
rect 1922 1731 1924 1733
rect 1932 1731 1942 1733
rect 1946 1731 1948 1733
rect 1956 1738 1958 1740
rect 1962 1738 1972 1740
rect 1980 1738 1982 1740
rect 1897 1715 1901 1723
rect 1935 1723 1939 1731
rect 1956 1730 1958 1732
rect 1962 1731 1965 1732
rect 1969 1731 1972 1732
rect 1962 1730 1972 1731
rect 1980 1730 1982 1732
rect 1888 1713 1890 1715
rect 1894 1713 1904 1715
rect 1912 1713 1914 1715
rect 1888 1705 1890 1707
rect 1894 1706 1897 1707
rect 1901 1706 1904 1707
rect 1894 1705 1904 1706
rect 1912 1705 1914 1707
rect 1922 1714 1924 1716
rect 1932 1715 1942 1716
rect 1932 1714 1935 1715
rect 1939 1714 1942 1715
rect 1946 1714 1948 1716
rect 1965 1715 1969 1723
rect 1922 1706 1924 1708
rect 1932 1706 1942 1708
rect 1946 1706 1948 1708
rect 1956 1713 1958 1715
rect 1962 1713 1972 1715
rect 1980 1713 1982 1715
rect 1897 1690 1901 1698
rect 1935 1698 1939 1706
rect 1956 1705 1958 1707
rect 1962 1706 1965 1707
rect 1969 1706 1972 1707
rect 1962 1705 1972 1706
rect 1980 1705 1982 1707
rect 1888 1688 1890 1690
rect 1894 1688 1904 1690
rect 1912 1688 1914 1690
rect 1888 1680 1890 1682
rect 1894 1681 1897 1682
rect 1901 1681 1904 1682
rect 1894 1680 1904 1681
rect 1912 1680 1914 1682
rect 1922 1689 1924 1691
rect 1932 1690 1942 1691
rect 1932 1689 1935 1690
rect 1939 1689 1942 1690
rect 1946 1689 1948 1691
rect 1965 1690 1969 1698
rect 1922 1681 1924 1683
rect 1932 1681 1942 1683
rect 1946 1681 1948 1683
rect 1956 1688 1958 1690
rect 1962 1688 1972 1690
rect 1980 1688 1982 1690
rect 1897 1665 1901 1673
rect 1935 1673 1939 1681
rect 1956 1680 1958 1682
rect 1962 1681 1965 1682
rect 1969 1681 1972 1682
rect 1962 1680 1972 1681
rect 1980 1680 1982 1682
rect 1888 1663 1890 1665
rect 1894 1663 1904 1665
rect 1912 1663 1914 1665
rect 1888 1655 1890 1657
rect 1894 1656 1897 1657
rect 1901 1656 1904 1657
rect 1894 1655 1904 1656
rect 1912 1655 1914 1657
rect 1922 1664 1924 1666
rect 1932 1665 1942 1666
rect 1932 1664 1935 1665
rect 1939 1664 1942 1665
rect 1946 1664 1948 1666
rect 1965 1665 1969 1673
rect 1922 1656 1924 1658
rect 1932 1656 1942 1658
rect 1946 1656 1948 1658
rect 1956 1663 1958 1665
rect 1962 1663 1972 1665
rect 1980 1663 1982 1665
rect 1897 1640 1901 1648
rect 1935 1648 1939 1656
rect 1956 1655 1958 1657
rect 1962 1656 1965 1657
rect 1969 1656 1972 1657
rect 1962 1655 1972 1656
rect 1980 1655 1982 1657
rect 1888 1638 1890 1640
rect 1894 1638 1904 1640
rect 1912 1638 1914 1640
rect 1888 1630 1890 1632
rect 1894 1631 1897 1632
rect 1901 1631 1904 1632
rect 1894 1630 1904 1631
rect 1912 1630 1914 1632
rect 1922 1639 1924 1641
rect 1932 1640 1942 1641
rect 1932 1639 1935 1640
rect 1939 1639 1942 1640
rect 1946 1639 1948 1641
rect 1965 1640 1969 1648
rect 1922 1631 1924 1633
rect 1932 1631 1942 1633
rect 1946 1631 1948 1633
rect 1956 1638 1958 1640
rect 1962 1638 1972 1640
rect 1980 1638 1982 1640
rect 1897 1615 1901 1623
rect 1935 1623 1939 1631
rect 1956 1630 1958 1632
rect 1962 1631 1965 1632
rect 1969 1631 1972 1632
rect 1962 1630 1972 1631
rect 1980 1630 1982 1632
rect 1888 1613 1890 1615
rect 1894 1613 1904 1615
rect 1912 1613 1914 1615
rect 1888 1605 1890 1607
rect 1894 1606 1897 1607
rect 1901 1606 1904 1607
rect 1894 1605 1904 1606
rect 1912 1605 1914 1607
rect 1922 1614 1924 1616
rect 1932 1615 1942 1616
rect 1932 1614 1935 1615
rect 1939 1614 1942 1615
rect 1946 1614 1948 1616
rect 1965 1615 1969 1623
rect 1922 1606 1924 1608
rect 1932 1606 1942 1608
rect 1946 1606 1948 1608
rect 1956 1613 1958 1615
rect 1962 1613 1972 1615
rect 1980 1613 1982 1615
rect 1897 1590 1901 1598
rect 1935 1598 1939 1606
rect 1956 1605 1958 1607
rect 1962 1606 1965 1607
rect 1969 1606 1972 1607
rect 1962 1605 1972 1606
rect 1980 1605 1982 1607
rect 1888 1588 1890 1590
rect 1894 1588 1904 1590
rect 1912 1588 1914 1590
rect 1888 1580 1890 1582
rect 1894 1581 1897 1582
rect 1901 1581 1904 1582
rect 1894 1580 1904 1581
rect 1912 1580 1914 1582
rect 1922 1589 1924 1591
rect 1932 1590 1942 1591
rect 1932 1589 1935 1590
rect 1939 1589 1942 1590
rect 1946 1589 1948 1591
rect 1965 1590 1969 1598
rect 1922 1581 1924 1583
rect 1932 1581 1942 1583
rect 1946 1581 1948 1583
rect 1956 1588 1958 1590
rect 1962 1588 1972 1590
rect 1980 1588 1982 1590
rect 1897 1565 1901 1573
rect 1935 1573 1939 1581
rect 1956 1580 1958 1582
rect 1962 1581 1965 1582
rect 1969 1581 1972 1582
rect 1962 1580 1972 1581
rect 1980 1580 1982 1582
rect 1888 1563 1890 1565
rect 1894 1563 1904 1565
rect 1912 1563 1914 1565
rect 1888 1555 1890 1557
rect 1894 1556 1897 1557
rect 1901 1556 1904 1557
rect 1894 1555 1904 1556
rect 1912 1555 1914 1557
rect 1922 1564 1924 1566
rect 1932 1565 1942 1566
rect 1932 1564 1935 1565
rect 1939 1564 1942 1565
rect 1946 1564 1948 1566
rect 1965 1565 1969 1573
rect 1922 1556 1924 1558
rect 1932 1556 1942 1558
rect 1946 1556 1948 1558
rect 1956 1563 1958 1565
rect 1962 1563 1972 1565
rect 1980 1563 1982 1565
rect 1897 1540 1901 1548
rect 1935 1548 1939 1556
rect 1956 1555 1958 1557
rect 1962 1556 1965 1557
rect 1969 1556 1972 1557
rect 1962 1555 1972 1556
rect 1980 1555 1982 1557
rect 1888 1538 1890 1540
rect 1894 1538 1904 1540
rect 1912 1538 1914 1540
rect 1888 1530 1890 1532
rect 1894 1531 1897 1532
rect 1901 1531 1904 1532
rect 1894 1530 1904 1531
rect 1912 1530 1914 1532
rect 1922 1539 1924 1541
rect 1932 1540 1942 1541
rect 1932 1539 1935 1540
rect 1939 1539 1942 1540
rect 1946 1539 1948 1541
rect 1965 1540 1969 1548
rect 1922 1531 1924 1533
rect 1932 1531 1942 1533
rect 1946 1531 1948 1533
rect 1956 1538 1958 1540
rect 1962 1538 1972 1540
rect 1980 1538 1982 1540
rect 1897 1515 1901 1523
rect 1935 1523 1939 1531
rect 1956 1530 1958 1532
rect 1962 1531 1965 1532
rect 1969 1531 1972 1532
rect 1962 1530 1972 1531
rect 1980 1530 1982 1532
rect 1888 1513 1890 1515
rect 1894 1513 1904 1515
rect 1912 1513 1914 1515
rect 1888 1505 1890 1507
rect 1894 1506 1897 1507
rect 1901 1506 1904 1507
rect 1894 1505 1904 1506
rect 1912 1505 1914 1507
rect 1922 1514 1924 1516
rect 1932 1515 1942 1516
rect 1932 1514 1935 1515
rect 1939 1514 1942 1515
rect 1946 1514 1948 1516
rect 1965 1515 1969 1523
rect 1922 1506 1924 1508
rect 1932 1506 1942 1508
rect 1946 1506 1948 1508
rect 1956 1513 1958 1515
rect 1962 1513 1972 1515
rect 1980 1513 1982 1515
rect 1897 1490 1901 1498
rect 1935 1498 1939 1506
rect 1956 1505 1958 1507
rect 1962 1506 1965 1507
rect 1969 1506 1972 1507
rect 1962 1505 1972 1506
rect 1980 1505 1982 1507
rect 1888 1488 1890 1490
rect 1894 1488 1904 1490
rect 1912 1488 1914 1490
rect 1888 1480 1890 1482
rect 1894 1481 1897 1482
rect 1901 1481 1904 1482
rect 1894 1480 1904 1481
rect 1912 1480 1914 1482
rect 1922 1489 1924 1491
rect 1932 1490 1942 1491
rect 1932 1489 1935 1490
rect 1939 1489 1942 1490
rect 1946 1489 1948 1491
rect 1965 1490 1969 1498
rect 1922 1481 1924 1483
rect 1932 1481 1942 1483
rect 1946 1481 1948 1483
rect 1956 1488 1958 1490
rect 1962 1488 1972 1490
rect 1980 1488 1982 1490
rect 1897 1465 1901 1473
rect 1935 1473 1939 1481
rect 1956 1480 1958 1482
rect 1962 1481 1965 1482
rect 1969 1481 1972 1482
rect 1962 1480 1972 1481
rect 1980 1480 1982 1482
rect 1888 1463 1890 1465
rect 1894 1463 1904 1465
rect 1912 1463 1914 1465
rect 1888 1455 1890 1457
rect 1894 1456 1897 1457
rect 1901 1456 1904 1457
rect 1894 1455 1904 1456
rect 1912 1455 1914 1457
rect 1922 1464 1924 1466
rect 1932 1465 1942 1466
rect 1932 1464 1935 1465
rect 1939 1464 1942 1465
rect 1946 1464 1948 1466
rect 1965 1465 1969 1473
rect 1922 1456 1924 1458
rect 1932 1456 1942 1458
rect 1946 1456 1948 1458
rect 1956 1463 1958 1465
rect 1962 1463 1972 1465
rect 1980 1463 1982 1465
rect 1897 1440 1901 1448
rect 1935 1448 1939 1456
rect 1956 1455 1958 1457
rect 1962 1456 1965 1457
rect 1969 1456 1972 1457
rect 1962 1455 1972 1456
rect 1980 1455 1982 1457
rect 1707 1433 1715 1434
rect 1710 1329 1712 1433
rect 1730 1410 1732 1434
rect 1740 1410 1742 1434
rect 1888 1438 1890 1440
rect 1894 1438 1904 1440
rect 1912 1438 1914 1440
rect 1888 1430 1890 1432
rect 1894 1431 1897 1432
rect 1901 1431 1904 1432
rect 1894 1430 1904 1431
rect 1912 1430 1914 1432
rect 1922 1439 1924 1441
rect 1932 1440 1942 1441
rect 1932 1439 1935 1440
rect 1939 1439 1942 1440
rect 1946 1439 1948 1441
rect 1965 1440 1969 1448
rect 1922 1431 1924 1433
rect 1932 1431 1942 1433
rect 1946 1431 1948 1433
rect 1956 1438 1958 1440
rect 1962 1438 1972 1440
rect 1980 1438 1982 1440
rect 1897 1415 1901 1423
rect 1935 1423 1939 1431
rect 1956 1430 1958 1432
rect 1962 1431 1965 1432
rect 1969 1431 1972 1432
rect 1962 1430 1972 1431
rect 1980 1430 1982 1432
rect 1758 1410 1760 1412
rect 1888 1413 1890 1415
rect 1894 1413 1904 1415
rect 1912 1413 1914 1415
rect 1888 1405 1890 1407
rect 1894 1406 1897 1407
rect 1901 1406 1904 1407
rect 1894 1405 1904 1406
rect 1912 1405 1914 1407
rect 1922 1414 1924 1416
rect 1932 1415 1942 1416
rect 1932 1414 1935 1415
rect 1939 1414 1942 1415
rect 1946 1414 1948 1416
rect 1965 1415 1969 1423
rect 1922 1406 1924 1408
rect 1932 1406 1942 1408
rect 1946 1406 1948 1408
rect 1956 1413 1958 1415
rect 1962 1413 1972 1415
rect 1980 1413 1982 1415
rect 1897 1390 1901 1398
rect 1935 1398 1939 1406
rect 1956 1405 1958 1407
rect 1962 1406 1965 1407
rect 1969 1406 1972 1407
rect 1962 1405 1972 1406
rect 1980 1405 1982 1407
rect 1758 1387 1760 1390
rect 1758 1383 1787 1387
rect 1758 1380 1760 1383
rect 1888 1388 1890 1390
rect 1894 1388 1904 1390
rect 1912 1388 1914 1390
rect 1888 1380 1890 1382
rect 1894 1381 1897 1382
rect 1901 1381 1904 1382
rect 1894 1380 1904 1381
rect 1912 1380 1914 1382
rect 1922 1389 1924 1391
rect 1932 1390 1942 1391
rect 1932 1389 1935 1390
rect 1939 1389 1942 1390
rect 1946 1389 1948 1391
rect 1965 1390 1969 1398
rect 1922 1381 1924 1383
rect 1932 1381 1942 1383
rect 1946 1381 1948 1383
rect 1956 1388 1958 1390
rect 1962 1388 1972 1390
rect 1980 1388 1982 1390
rect 1758 1368 1760 1370
rect 1897 1365 1901 1373
rect 1935 1373 1939 1381
rect 1956 1380 1958 1382
rect 1962 1381 1965 1382
rect 1969 1381 1972 1382
rect 1962 1380 1972 1381
rect 1980 1380 1982 1382
rect 1730 1328 1732 1365
rect 1740 1329 1742 1362
rect 1888 1363 1890 1365
rect 1894 1363 1904 1365
rect 1912 1363 1914 1365
rect 1888 1355 1890 1357
rect 1894 1356 1897 1357
rect 1901 1356 1904 1357
rect 1894 1355 1904 1356
rect 1912 1355 1914 1357
rect 1922 1364 1924 1366
rect 1932 1365 1942 1366
rect 1932 1364 1935 1365
rect 1939 1364 1942 1365
rect 1946 1364 1948 1366
rect 1965 1365 1969 1373
rect 1922 1356 1924 1358
rect 1932 1356 1942 1358
rect 1946 1356 1948 1358
rect 1956 1363 1958 1365
rect 1962 1363 1972 1365
rect 1980 1363 1982 1365
rect 1897 1340 1901 1348
rect 1935 1348 1939 1356
rect 1956 1355 1958 1357
rect 1962 1356 1965 1357
rect 1969 1356 1972 1357
rect 1962 1355 1972 1356
rect 1980 1355 1982 1357
rect 1888 1338 1890 1340
rect 1894 1338 1904 1340
rect 1912 1338 1914 1340
rect 1888 1330 1890 1332
rect 1894 1331 1897 1332
rect 1901 1331 1904 1332
rect 1894 1330 1904 1331
rect 1912 1330 1914 1332
rect 1922 1339 1924 1341
rect 1932 1340 1942 1341
rect 1932 1339 1935 1340
rect 1939 1339 1942 1340
rect 1946 1339 1948 1341
rect 1965 1340 1969 1348
rect 1922 1331 1924 1333
rect 1932 1331 1942 1333
rect 1946 1331 1948 1333
rect 1956 1338 1958 1340
rect 1962 1338 1972 1340
rect 1980 1338 1982 1340
rect 1897 1315 1901 1323
rect 1935 1323 1939 1331
rect 1956 1330 1958 1332
rect 1962 1331 1965 1332
rect 1969 1331 1972 1332
rect 1962 1330 1972 1331
rect 1980 1330 1982 1332
rect 1888 1313 1890 1315
rect 1894 1313 1904 1315
rect 1912 1313 1914 1315
rect 1888 1305 1890 1307
rect 1894 1306 1897 1307
rect 1901 1306 1904 1307
rect 1894 1305 1904 1306
rect 1912 1305 1914 1307
rect 1922 1314 1924 1316
rect 1932 1315 1942 1316
rect 1932 1314 1935 1315
rect 1939 1314 1942 1315
rect 1946 1314 1948 1316
rect 1965 1315 1969 1323
rect 1922 1306 1924 1308
rect 1932 1306 1942 1308
rect 1946 1306 1948 1308
rect 1956 1313 1958 1315
rect 1962 1313 1972 1315
rect 1980 1313 1982 1315
rect 1897 1290 1901 1298
rect 1935 1298 1939 1306
rect 1956 1305 1958 1307
rect 1962 1306 1965 1307
rect 1969 1306 1972 1307
rect 1962 1305 1972 1306
rect 1980 1305 1982 1307
rect 1888 1288 1890 1290
rect 1894 1288 1904 1290
rect 1912 1288 1914 1290
rect 1888 1280 1890 1282
rect 1894 1281 1897 1282
rect 1901 1281 1904 1282
rect 1894 1280 1904 1281
rect 1912 1280 1914 1282
rect 1922 1289 1924 1291
rect 1932 1290 1942 1291
rect 1932 1289 1935 1290
rect 1939 1289 1942 1290
rect 1946 1289 1948 1291
rect 1965 1290 1969 1298
rect 1922 1281 1924 1283
rect 1932 1281 1942 1283
rect 1946 1281 1948 1283
rect 1956 1288 1958 1290
rect 1962 1288 1972 1290
rect 1980 1288 1982 1290
rect 1897 1265 1901 1273
rect 1935 1273 1939 1281
rect 1956 1280 1958 1282
rect 1962 1281 1965 1282
rect 1969 1281 1972 1282
rect 1962 1280 1972 1281
rect 1980 1280 1982 1282
rect 1888 1263 1890 1265
rect 1894 1263 1904 1265
rect 1912 1263 1914 1265
rect 1888 1255 1890 1257
rect 1894 1256 1897 1257
rect 1901 1256 1904 1257
rect 1894 1255 1904 1256
rect 1912 1255 1914 1257
rect 1922 1264 1924 1266
rect 1932 1265 1942 1266
rect 1932 1264 1935 1265
rect 1939 1264 1942 1265
rect 1946 1264 1948 1266
rect 1965 1265 1969 1273
rect 1922 1256 1924 1258
rect 1932 1256 1942 1258
rect 1946 1256 1948 1258
rect 1956 1263 1958 1265
rect 1962 1263 1972 1265
rect 1980 1263 1982 1265
rect 1897 1240 1901 1248
rect 1935 1248 1939 1256
rect 1956 1255 1958 1257
rect 1962 1256 1965 1257
rect 1969 1256 1972 1257
rect 1962 1255 1972 1256
rect 1980 1255 1982 1257
rect 1888 1238 1890 1240
rect 1894 1238 1904 1240
rect 1912 1238 1914 1240
rect 1888 1230 1890 1232
rect 1894 1231 1897 1232
rect 1901 1231 1904 1232
rect 1894 1230 1904 1231
rect 1912 1230 1914 1232
rect 1922 1239 1924 1241
rect 1932 1240 1942 1241
rect 1932 1239 1935 1240
rect 1939 1239 1942 1240
rect 1946 1239 1948 1241
rect 1965 1240 1969 1248
rect 1922 1231 1924 1233
rect 1932 1231 1942 1233
rect 1946 1231 1948 1233
rect 1956 1238 1958 1240
rect 1962 1238 1972 1240
rect 1980 1238 1982 1240
rect 1897 1215 1901 1223
rect 1935 1223 1939 1231
rect 1956 1230 1958 1232
rect 1962 1231 1965 1232
rect 1969 1231 1972 1232
rect 1962 1230 1972 1231
rect 1980 1230 1982 1232
rect 1888 1213 1890 1215
rect 1894 1213 1904 1215
rect 1912 1213 1914 1215
rect 1888 1205 1890 1207
rect 1894 1206 1897 1207
rect 1901 1206 1904 1207
rect 1894 1205 1904 1206
rect 1912 1205 1914 1207
rect 1922 1214 1924 1216
rect 1932 1215 1942 1216
rect 1932 1214 1935 1215
rect 1939 1214 1942 1215
rect 1946 1214 1948 1216
rect 1965 1215 1969 1223
rect 1922 1206 1924 1208
rect 1932 1206 1942 1208
rect 1946 1206 1948 1208
rect 1956 1213 1958 1215
rect 1962 1213 1972 1215
rect 1980 1213 1982 1215
rect 912 1198 914 1200
rect 1897 1190 1901 1198
rect 1935 1198 1939 1206
rect 1956 1205 1958 1207
rect 1962 1206 1965 1207
rect 1969 1206 1972 1207
rect 1962 1205 1972 1206
rect 1980 1205 1982 1207
rect 912 1178 914 1188
rect 1888 1188 1890 1190
rect 1894 1188 1904 1190
rect 1912 1188 1914 1190
rect 1888 1180 1890 1182
rect 1894 1181 1897 1182
rect 1901 1181 1904 1182
rect 1894 1180 1904 1181
rect 1912 1180 1914 1182
rect 1922 1189 1924 1191
rect 1932 1190 1942 1191
rect 1932 1189 1935 1190
rect 1939 1189 1942 1190
rect 1946 1189 1948 1191
rect 1965 1190 1969 1198
rect 1922 1181 1924 1183
rect 1932 1181 1942 1183
rect 1946 1181 1948 1183
rect 1956 1188 1958 1190
rect 1962 1188 1972 1190
rect 1980 1188 1982 1190
rect 1897 1165 1901 1173
rect 1935 1173 1939 1181
rect 1956 1180 1958 1182
rect 1962 1181 1965 1182
rect 1969 1181 1972 1182
rect 1962 1180 1972 1181
rect 1980 1180 1982 1182
rect 912 1156 914 1158
rect 1888 1163 1890 1165
rect 1894 1163 1904 1165
rect 1912 1163 1914 1165
rect 1888 1155 1890 1157
rect 1894 1156 1897 1157
rect 1901 1156 1904 1157
rect 1894 1155 1904 1156
rect 1912 1155 1914 1157
rect 1922 1164 1924 1166
rect 1932 1165 1942 1166
rect 1932 1164 1935 1165
rect 1939 1164 1942 1165
rect 1946 1164 1948 1166
rect 1965 1165 1969 1173
rect 1922 1156 1924 1158
rect 1932 1156 1942 1158
rect 1946 1156 1948 1158
rect 1956 1163 1958 1165
rect 1962 1163 1972 1165
rect 1980 1163 1982 1165
rect 1897 1140 1901 1148
rect 1935 1148 1939 1156
rect 1956 1155 1958 1157
rect 1962 1156 1965 1157
rect 1969 1156 1972 1157
rect 1962 1155 1972 1156
rect 1980 1155 1982 1157
rect 1888 1138 1890 1140
rect 1894 1138 1904 1140
rect 1912 1138 1914 1140
rect 1888 1130 1890 1132
rect 1894 1131 1897 1132
rect 1901 1131 1904 1132
rect 1894 1130 1904 1131
rect 1912 1130 1914 1132
rect 1922 1139 1924 1141
rect 1932 1140 1942 1141
rect 1932 1139 1935 1140
rect 1939 1139 1942 1140
rect 1946 1139 1948 1141
rect 1965 1140 1969 1148
rect 1922 1131 1924 1133
rect 1932 1131 1942 1133
rect 1946 1131 1948 1133
rect 1956 1138 1958 1140
rect 1962 1138 1972 1140
rect 1980 1138 1982 1140
rect 1897 1115 1901 1123
rect 1935 1123 1939 1131
rect 1956 1130 1958 1132
rect 1962 1131 1965 1132
rect 1969 1131 1972 1132
rect 1962 1130 1972 1131
rect 1980 1130 1982 1132
rect 1888 1113 1890 1115
rect 1894 1113 1904 1115
rect 1912 1113 1914 1115
rect 1888 1105 1890 1107
rect 1894 1106 1897 1107
rect 1901 1106 1904 1107
rect 1894 1105 1904 1106
rect 1912 1105 1914 1107
rect 1922 1114 1924 1116
rect 1932 1115 1942 1116
rect 1932 1114 1935 1115
rect 1939 1114 1942 1115
rect 1946 1114 1948 1116
rect 1965 1115 1969 1123
rect 1922 1106 1924 1108
rect 1932 1106 1942 1108
rect 1946 1106 1948 1108
rect 1956 1113 1958 1115
rect 1962 1113 1972 1115
rect 1980 1113 1982 1115
rect 1754 1097 1755 1101
rect 1735 1093 1737 1095
rect 1753 1093 1755 1097
rect 1763 1097 1764 1101
rect 1763 1093 1765 1097
rect 1897 1090 1901 1098
rect 1935 1098 1939 1106
rect 1956 1105 1958 1107
rect 1962 1106 1965 1107
rect 1969 1106 1972 1107
rect 1962 1105 1972 1106
rect 1980 1105 1982 1107
rect 1888 1088 1890 1090
rect 1894 1088 1904 1090
rect 1912 1088 1914 1090
rect 1888 1080 1890 1082
rect 1894 1081 1897 1082
rect 1901 1081 1904 1082
rect 1894 1080 1904 1081
rect 1912 1080 1914 1082
rect 1922 1089 1924 1091
rect 1932 1090 1942 1091
rect 1932 1089 1935 1090
rect 1939 1089 1942 1090
rect 1946 1089 1948 1091
rect 1965 1090 1969 1098
rect 1922 1081 1924 1083
rect 1932 1081 1942 1083
rect 1946 1081 1948 1083
rect 1956 1088 1958 1090
rect 1962 1088 1972 1090
rect 1980 1088 1982 1090
rect 1735 1072 1737 1075
rect 1735 1068 1736 1072
rect 1735 1065 1737 1068
rect 1753 1065 1755 1075
rect 1763 1065 1765 1075
rect 1897 1065 1901 1073
rect 1935 1073 1939 1081
rect 1956 1080 1958 1082
rect 1962 1081 1965 1082
rect 1969 1081 1972 1082
rect 1962 1080 1972 1081
rect 1980 1080 1982 1082
rect 1888 1063 1890 1065
rect 1894 1063 1904 1065
rect 1912 1063 1914 1065
rect 1888 1055 1890 1057
rect 1894 1056 1897 1057
rect 1901 1056 1904 1057
rect 1894 1055 1904 1056
rect 1912 1055 1914 1057
rect 1922 1064 1924 1066
rect 1932 1065 1942 1066
rect 1932 1064 1935 1065
rect 1939 1064 1942 1065
rect 1946 1064 1948 1066
rect 1965 1065 1969 1073
rect 1922 1056 1924 1058
rect 1932 1056 1942 1058
rect 1946 1056 1948 1058
rect 1956 1063 1958 1065
rect 1962 1063 1972 1065
rect 1980 1063 1982 1065
rect 1735 1053 1737 1055
rect 1753 1053 1755 1055
rect 1763 1053 1765 1055
rect 1897 1040 1901 1048
rect 1935 1048 1939 1056
rect 1956 1055 1958 1057
rect 1962 1056 1965 1057
rect 1969 1056 1972 1057
rect 1962 1055 1972 1056
rect 1980 1055 1982 1057
rect 1888 1038 1890 1040
rect 1894 1038 1904 1040
rect 1912 1038 1914 1040
rect 1888 1030 1890 1032
rect 1894 1031 1897 1032
rect 1901 1031 1904 1032
rect 1894 1030 1904 1031
rect 1912 1030 1914 1032
rect 1922 1039 1924 1041
rect 1932 1040 1942 1041
rect 1932 1039 1935 1040
rect 1939 1039 1942 1040
rect 1946 1039 1948 1041
rect 1965 1040 1969 1048
rect 1922 1031 1924 1033
rect 1932 1031 1942 1033
rect 1946 1031 1948 1033
rect 1956 1038 1958 1040
rect 1962 1038 1972 1040
rect 1980 1038 1982 1040
rect 1897 1015 1901 1023
rect 1935 1023 1939 1031
rect 1956 1030 1958 1032
rect 1962 1031 1965 1032
rect 1969 1031 1972 1032
rect 1962 1030 1972 1031
rect 1980 1030 1982 1032
rect 1888 1013 1890 1015
rect 1894 1013 1904 1015
rect 1912 1013 1914 1015
rect 1888 1005 1890 1007
rect 1894 1006 1897 1007
rect 1901 1006 1904 1007
rect 1894 1005 1904 1006
rect 1912 1005 1914 1007
rect 1922 1014 1924 1016
rect 1932 1015 1942 1016
rect 1932 1014 1935 1015
rect 1939 1014 1942 1015
rect 1946 1014 1948 1016
rect 1965 1015 1969 1023
rect 1922 1006 1924 1008
rect 1932 1006 1942 1008
rect 1946 1006 1948 1008
rect 1956 1013 1958 1015
rect 1962 1013 1972 1015
rect 1980 1013 1982 1015
rect 1897 990 1901 998
rect 1935 998 1939 1006
rect 1956 1005 1958 1007
rect 1962 1006 1965 1007
rect 1969 1006 1972 1007
rect 1962 1005 1972 1006
rect 1980 1005 1982 1007
rect 1888 988 1890 990
rect 1894 988 1904 990
rect 1912 988 1914 990
rect 1888 980 1890 982
rect 1894 981 1897 982
rect 1901 981 1904 982
rect 1894 980 1904 981
rect 1912 980 1914 982
rect 1922 989 1924 991
rect 1932 990 1942 991
rect 1932 989 1935 990
rect 1939 989 1942 990
rect 1946 989 1948 991
rect 1965 990 1969 998
rect 1922 981 1924 983
rect 1932 981 1942 983
rect 1946 981 1948 983
rect 1956 988 1958 990
rect 1962 988 1972 990
rect 1980 988 1982 990
rect 1897 965 1901 973
rect 1935 973 1939 981
rect 1956 980 1958 982
rect 1962 981 1965 982
rect 1969 981 1972 982
rect 1962 980 1972 981
rect 1980 980 1982 982
rect 1888 963 1890 965
rect 1894 963 1904 965
rect 1912 963 1914 965
rect 1888 955 1890 957
rect 1894 956 1897 957
rect 1901 956 1904 957
rect 1894 955 1904 956
rect 1912 955 1914 957
rect 1922 964 1924 966
rect 1932 965 1942 966
rect 1932 964 1935 965
rect 1939 964 1942 965
rect 1946 964 1948 966
rect 1965 965 1969 973
rect 1922 956 1924 958
rect 1932 956 1942 958
rect 1946 956 1948 958
rect 1956 963 1958 965
rect 1962 963 1972 965
rect 1980 963 1982 965
rect 1897 940 1901 948
rect 1935 948 1939 956
rect 1956 955 1958 957
rect 1962 956 1965 957
rect 1969 956 1972 957
rect 1962 955 1972 956
rect 1980 955 1982 957
rect 1888 938 1890 940
rect 1894 938 1904 940
rect 1912 938 1914 940
rect 1888 930 1890 932
rect 1894 931 1897 932
rect 1901 931 1904 932
rect 1894 930 1904 931
rect 1912 930 1914 932
rect 1922 939 1924 941
rect 1932 940 1942 941
rect 1932 939 1935 940
rect 1939 939 1942 940
rect 1946 939 1948 941
rect 1965 940 1969 948
rect 1922 931 1924 933
rect 1932 931 1942 933
rect 1946 931 1948 933
rect 1956 938 1958 940
rect 1962 938 1972 940
rect 1980 938 1982 940
rect 1897 915 1901 923
rect 1935 923 1939 931
rect 1956 930 1958 932
rect 1962 931 1965 932
rect 1969 931 1972 932
rect 1962 930 1972 931
rect 1980 930 1982 932
rect 1888 913 1890 915
rect 1894 913 1904 915
rect 1912 913 1914 915
rect 1888 905 1890 907
rect 1894 906 1897 907
rect 1901 906 1904 907
rect 1894 905 1904 906
rect 1912 905 1914 907
rect 1922 914 1924 916
rect 1932 915 1942 916
rect 1932 914 1935 915
rect 1939 914 1942 915
rect 1946 914 1948 916
rect 1965 915 1969 923
rect 1922 906 1924 908
rect 1932 906 1942 908
rect 1946 906 1948 908
rect 1956 913 1958 915
rect 1962 913 1972 915
rect 1980 913 1982 915
rect 1897 890 1901 898
rect 1935 898 1939 906
rect 1956 905 1958 907
rect 1962 906 1965 907
rect 1969 906 1972 907
rect 1962 905 1972 906
rect 1980 905 1982 907
rect 1888 888 1890 890
rect 1894 888 1904 890
rect 1912 888 1914 890
rect 1888 880 1890 882
rect 1894 881 1897 882
rect 1901 881 1904 882
rect 1894 880 1904 881
rect 1912 880 1914 882
rect 1922 889 1924 891
rect 1932 890 1942 891
rect 1932 889 1935 890
rect 1939 889 1942 890
rect 1946 889 1948 891
rect 1965 890 1969 898
rect 1922 881 1924 883
rect 1932 881 1942 883
rect 1946 881 1948 883
rect 1956 888 1958 890
rect 1962 888 1972 890
rect 1980 888 1982 890
rect 1897 865 1901 873
rect 1935 873 1939 881
rect 1956 880 1958 882
rect 1962 881 1965 882
rect 1969 881 1972 882
rect 1962 880 1972 881
rect 1980 880 1982 882
rect 1888 863 1890 865
rect 1894 863 1904 865
rect 1912 863 1914 865
rect 1888 855 1890 857
rect 1894 856 1897 857
rect 1901 856 1904 857
rect 1894 855 1904 856
rect 1912 855 1914 857
rect 1922 864 1924 866
rect 1932 865 1942 866
rect 1932 864 1935 865
rect 1939 864 1942 865
rect 1946 864 1948 866
rect 1965 865 1969 873
rect 1922 856 1924 858
rect 1932 856 1942 858
rect 1946 856 1948 858
rect 1956 863 1958 865
rect 1962 863 1972 865
rect 1980 863 1982 865
rect 1897 840 1901 848
rect 1935 848 1939 856
rect 1956 855 1958 857
rect 1962 856 1965 857
rect 1969 856 1972 857
rect 1962 855 1972 856
rect 1980 855 1982 857
rect 1888 838 1890 840
rect 1894 838 1904 840
rect 1912 838 1914 840
rect 1888 830 1890 832
rect 1894 831 1897 832
rect 1901 831 1904 832
rect 1894 830 1904 831
rect 1912 830 1914 832
rect 1922 839 1924 841
rect 1932 840 1942 841
rect 1932 839 1935 840
rect 1939 839 1942 840
rect 1946 839 1948 841
rect 1965 840 1969 848
rect 1922 831 1924 833
rect 1932 831 1942 833
rect 1946 831 1948 833
rect 1956 838 1958 840
rect 1962 838 1972 840
rect 1980 838 1982 840
rect 1897 815 1901 823
rect 1935 823 1939 831
rect 1956 830 1958 832
rect 1962 831 1965 832
rect 1969 831 1972 832
rect 1962 830 1972 831
rect 1980 830 1982 832
rect 1888 813 1890 815
rect 1894 813 1904 815
rect 1912 813 1914 815
rect 1888 805 1890 807
rect 1894 806 1897 807
rect 1901 806 1904 807
rect 1894 805 1904 806
rect 1912 805 1914 807
rect 1922 814 1924 816
rect 1932 815 1942 816
rect 1932 814 1935 815
rect 1939 814 1942 815
rect 1946 814 1948 816
rect 1965 815 1969 823
rect 1922 806 1924 808
rect 1932 806 1942 808
rect 1946 806 1948 808
rect 1956 813 1958 815
rect 1962 813 1972 815
rect 1980 813 1982 815
rect 1897 790 1901 798
rect 1935 798 1939 806
rect 1956 805 1958 807
rect 1962 806 1965 807
rect 1969 806 1972 807
rect 1962 805 1972 806
rect 1980 805 1982 807
rect 1888 788 1890 790
rect 1894 788 1904 790
rect 1912 788 1914 790
rect 1888 780 1890 782
rect 1894 781 1897 782
rect 1901 781 1904 782
rect 1894 780 1904 781
rect 1912 780 1914 782
rect 1922 789 1924 791
rect 1932 790 1942 791
rect 1932 789 1935 790
rect 1939 789 1942 790
rect 1946 789 1948 791
rect 1965 790 1969 798
rect 1922 781 1924 783
rect 1932 781 1942 783
rect 1946 781 1948 783
rect 1956 788 1958 790
rect 1962 788 1972 790
rect 1980 788 1982 790
rect 1897 765 1901 773
rect 1935 773 1939 781
rect 1956 780 1958 782
rect 1962 781 1965 782
rect 1969 781 1972 782
rect 1962 780 1972 781
rect 1980 780 1982 782
rect 1888 763 1890 765
rect 1894 763 1904 765
rect 1912 763 1914 765
rect 1888 755 1890 757
rect 1894 756 1897 757
rect 1901 756 1904 757
rect 1894 755 1904 756
rect 1912 755 1914 757
rect 1922 764 1924 766
rect 1932 765 1942 766
rect 1932 764 1935 765
rect 1939 764 1942 765
rect 1946 764 1948 766
rect 1965 765 1969 773
rect 1922 756 1924 758
rect 1932 756 1942 758
rect 1946 756 1948 758
rect 1956 763 1958 765
rect 1962 763 1972 765
rect 1980 763 1982 765
rect 1897 740 1901 748
rect 1935 748 1939 756
rect 1956 755 1958 757
rect 1962 756 1965 757
rect 1969 756 1972 757
rect 1962 755 1972 756
rect 1980 755 1982 757
rect 1888 738 1890 740
rect 1894 738 1904 740
rect 1912 738 1914 740
rect 1888 730 1890 732
rect 1894 731 1897 732
rect 1901 731 1904 732
rect 1894 730 1904 731
rect 1912 730 1914 732
rect 1922 739 1924 741
rect 1932 740 1942 741
rect 1932 739 1935 740
rect 1939 739 1942 740
rect 1946 739 1948 741
rect 1965 740 1969 748
rect 1922 731 1924 733
rect 1932 731 1942 733
rect 1946 731 1948 733
rect 1956 738 1958 740
rect 1962 738 1972 740
rect 1980 738 1982 740
rect 1897 715 1901 723
rect 1935 723 1939 731
rect 1956 730 1958 732
rect 1962 731 1965 732
rect 1969 731 1972 732
rect 1962 730 1972 731
rect 1980 730 1982 732
rect 1888 713 1890 715
rect 1894 713 1904 715
rect 1912 713 1914 715
rect 1888 705 1890 707
rect 1894 706 1897 707
rect 1901 706 1904 707
rect 1894 705 1904 706
rect 1912 705 1914 707
rect 1922 714 1924 716
rect 1932 715 1942 716
rect 1932 714 1935 715
rect 1939 714 1942 715
rect 1946 714 1948 716
rect 1965 715 1969 723
rect 1922 706 1924 708
rect 1932 706 1942 708
rect 1946 706 1948 708
rect 1956 713 1958 715
rect 1962 713 1972 715
rect 1980 713 1982 715
rect 1897 690 1901 698
rect 1935 698 1939 706
rect 1956 705 1958 707
rect 1962 706 1965 707
rect 1969 706 1972 707
rect 1962 705 1972 706
rect 1980 705 1982 707
rect 1888 688 1890 690
rect 1894 688 1904 690
rect 1912 688 1914 690
rect 1888 680 1890 682
rect 1894 681 1897 682
rect 1901 681 1904 682
rect 1894 680 1904 681
rect 1912 680 1914 682
rect 1922 689 1924 691
rect 1932 690 1942 691
rect 1932 689 1935 690
rect 1939 689 1942 690
rect 1946 689 1948 691
rect 1965 690 1969 698
rect 1922 681 1924 683
rect 1932 681 1942 683
rect 1946 681 1948 683
rect 1956 688 1958 690
rect 1962 688 1972 690
rect 1980 688 1982 690
rect 1897 665 1901 673
rect 1935 673 1939 681
rect 1956 680 1958 682
rect 1962 681 1965 682
rect 1969 681 1972 682
rect 1962 680 1972 681
rect 1980 680 1982 682
rect 1888 663 1890 665
rect 1894 663 1904 665
rect 1912 663 1914 665
rect 1888 655 1890 657
rect 1894 656 1897 657
rect 1901 656 1904 657
rect 1894 655 1904 656
rect 1912 655 1914 657
rect 1922 664 1924 666
rect 1932 665 1942 666
rect 1932 664 1935 665
rect 1939 664 1942 665
rect 1946 664 1948 666
rect 1965 665 1969 673
rect 1922 656 1924 658
rect 1932 656 1942 658
rect 1946 656 1948 658
rect 1956 663 1958 665
rect 1962 663 1972 665
rect 1980 663 1982 665
rect 1897 640 1901 648
rect 1935 648 1939 656
rect 1956 655 1958 657
rect 1962 656 1965 657
rect 1969 656 1972 657
rect 1962 655 1972 656
rect 1980 655 1982 657
rect 1888 638 1890 640
rect 1894 638 1904 640
rect 1912 638 1914 640
rect 1888 630 1890 632
rect 1894 631 1897 632
rect 1901 631 1904 632
rect 1894 630 1904 631
rect 1912 630 1914 632
rect 1922 639 1924 641
rect 1932 640 1942 641
rect 1932 639 1935 640
rect 1939 639 1942 640
rect 1946 639 1948 641
rect 1965 640 1969 648
rect 1922 631 1924 633
rect 1932 631 1942 633
rect 1946 631 1948 633
rect 1956 638 1958 640
rect 1962 638 1972 640
rect 1980 638 1982 640
rect 1897 615 1901 623
rect 1935 623 1939 631
rect 1956 630 1958 632
rect 1962 631 1965 632
rect 1969 631 1972 632
rect 1962 630 1972 631
rect 1980 630 1982 632
rect 1888 613 1890 615
rect 1894 613 1904 615
rect 1912 613 1914 615
rect 1888 605 1890 607
rect 1894 606 1897 607
rect 1901 606 1904 607
rect 1894 605 1904 606
rect 1912 605 1914 607
rect 1922 614 1924 616
rect 1932 615 1942 616
rect 1932 614 1935 615
rect 1939 614 1942 615
rect 1946 614 1948 616
rect 1965 615 1969 623
rect 1922 606 1924 608
rect 1932 606 1942 608
rect 1946 606 1948 608
rect 1956 613 1958 615
rect 1962 613 1972 615
rect 1980 613 1982 615
rect 1897 590 1901 598
rect 1935 598 1939 606
rect 1956 605 1958 607
rect 1962 606 1965 607
rect 1969 606 1972 607
rect 1962 605 1972 606
rect 1980 605 1982 607
rect 1888 588 1890 590
rect 1894 588 1904 590
rect 1912 588 1914 590
rect 1888 580 1890 582
rect 1894 581 1897 582
rect 1901 581 1904 582
rect 1894 580 1904 581
rect 1912 580 1914 582
rect 1922 589 1924 591
rect 1932 590 1942 591
rect 1932 589 1935 590
rect 1939 589 1942 590
rect 1946 589 1948 591
rect 1965 590 1969 598
rect 1922 581 1924 583
rect 1932 581 1942 583
rect 1946 581 1948 583
rect 1956 588 1958 590
rect 1962 588 1972 590
rect 1980 588 1982 590
rect 1897 565 1901 573
rect 1935 573 1939 581
rect 1956 580 1958 582
rect 1962 581 1965 582
rect 1969 581 1972 582
rect 1962 580 1972 581
rect 1980 580 1982 582
rect 1888 563 1890 565
rect 1894 563 1904 565
rect 1912 563 1914 565
rect 1888 555 1890 557
rect 1894 556 1897 557
rect 1901 556 1904 557
rect 1894 555 1904 556
rect 1912 555 1914 557
rect 1922 564 1924 566
rect 1932 565 1942 566
rect 1932 564 1935 565
rect 1939 564 1942 565
rect 1946 564 1948 566
rect 1965 565 1969 573
rect 1922 556 1924 558
rect 1932 556 1942 558
rect 1946 556 1948 558
rect 1956 563 1958 565
rect 1962 563 1972 565
rect 1980 563 1982 565
rect 1897 540 1901 548
rect 1935 548 1939 556
rect 1956 555 1958 557
rect 1962 556 1965 557
rect 1969 556 1972 557
rect 1962 555 1972 556
rect 1980 555 1982 557
rect 1888 538 1890 540
rect 1894 538 1904 540
rect 1912 538 1914 540
rect 1888 530 1890 532
rect 1894 531 1897 532
rect 1901 531 1904 532
rect 1894 530 1904 531
rect 1912 530 1914 532
rect 1922 539 1924 541
rect 1932 540 1942 541
rect 1932 539 1935 540
rect 1939 539 1942 540
rect 1946 539 1948 541
rect 1965 540 1969 548
rect 1922 531 1924 533
rect 1932 531 1942 533
rect 1946 531 1948 533
rect 1956 538 1958 540
rect 1962 538 1972 540
rect 1980 538 1982 540
rect 1897 515 1901 523
rect 1935 523 1939 531
rect 1956 530 1958 532
rect 1962 531 1965 532
rect 1969 531 1972 532
rect 1962 530 1972 531
rect 1980 530 1982 532
rect 1888 513 1890 515
rect 1894 513 1904 515
rect 1912 513 1914 515
rect 1888 505 1890 507
rect 1894 506 1897 507
rect 1901 506 1904 507
rect 1894 505 1904 506
rect 1912 505 1914 507
rect 1922 514 1924 516
rect 1932 515 1942 516
rect 1932 514 1935 515
rect 1939 514 1942 515
rect 1946 514 1948 516
rect 1965 515 1969 523
rect 1922 506 1924 508
rect 1932 506 1942 508
rect 1946 506 1948 508
rect 1956 513 1958 515
rect 1962 513 1972 515
rect 1980 513 1982 515
rect 1897 490 1901 498
rect 1935 498 1939 506
rect 1956 505 1958 507
rect 1962 506 1965 507
rect 1969 506 1972 507
rect 1962 505 1972 506
rect 1980 505 1982 507
rect 1888 488 1890 490
rect 1894 488 1904 490
rect 1912 488 1914 490
rect 1888 480 1890 482
rect 1894 481 1897 482
rect 1901 481 1904 482
rect 1894 480 1904 481
rect 1912 480 1914 482
rect 1922 489 1924 491
rect 1932 490 1942 491
rect 1932 489 1935 490
rect 1939 489 1942 490
rect 1946 489 1948 491
rect 1965 490 1969 498
rect 1922 481 1924 483
rect 1932 481 1942 483
rect 1946 481 1948 483
rect 1956 488 1958 490
rect 1962 488 1972 490
rect 1980 488 1982 490
rect 1897 465 1901 473
rect 1935 473 1939 481
rect 1956 480 1958 482
rect 1962 481 1965 482
rect 1969 481 1972 482
rect 1962 480 1972 481
rect 1980 480 1982 482
rect 1888 463 1890 465
rect 1894 463 1904 465
rect 1912 463 1914 465
rect 1888 455 1890 457
rect 1894 456 1897 457
rect 1901 456 1904 457
rect 1894 455 1904 456
rect 1912 455 1914 457
rect 1922 464 1924 466
rect 1932 465 1942 466
rect 1932 464 1935 465
rect 1939 464 1942 465
rect 1946 464 1948 466
rect 1965 465 1969 473
rect 1922 456 1924 458
rect 1932 456 1942 458
rect 1946 456 1948 458
rect 1956 463 1958 465
rect 1962 463 1972 465
rect 1980 463 1982 465
rect 1897 440 1901 448
rect 1935 448 1939 456
rect 1956 455 1958 457
rect 1962 456 1965 457
rect 1969 456 1972 457
rect 1962 455 1972 456
rect 1980 455 1982 457
rect 1888 438 1890 440
rect 1894 438 1904 440
rect 1912 438 1914 440
rect 1888 430 1890 432
rect 1894 431 1897 432
rect 1901 431 1904 432
rect 1894 430 1904 431
rect 1912 430 1914 432
rect 1922 439 1924 441
rect 1932 440 1942 441
rect 1932 439 1935 440
rect 1939 439 1942 440
rect 1946 439 1948 441
rect 1965 440 1969 448
rect 1922 431 1924 433
rect 1932 431 1942 433
rect 1946 431 1948 433
rect 1956 438 1958 440
rect 1962 438 1972 440
rect 1980 438 1982 440
rect 1897 415 1901 423
rect 1935 423 1939 431
rect 1956 430 1958 432
rect 1962 431 1965 432
rect 1969 431 1972 432
rect 1962 430 1972 431
rect 1980 430 1982 432
rect 1888 413 1890 415
rect 1894 413 1904 415
rect 1912 413 1914 415
rect 1888 405 1890 407
rect 1894 406 1897 407
rect 1901 406 1904 407
rect 1894 405 1904 406
rect 1912 405 1914 407
rect 1922 414 1924 416
rect 1932 415 1942 416
rect 1932 414 1935 415
rect 1939 414 1942 415
rect 1946 414 1948 416
rect 1965 415 1969 423
rect 1922 406 1924 408
rect 1932 406 1942 408
rect 1946 406 1948 408
rect 1956 413 1958 415
rect 1962 413 1972 415
rect 1980 413 1982 415
rect 1897 390 1901 398
rect 1935 398 1939 406
rect 1956 405 1958 407
rect 1962 406 1965 407
rect 1969 406 1972 407
rect 1962 405 1972 406
rect 1980 405 1982 407
rect 1888 388 1890 390
rect 1894 388 1904 390
rect 1912 388 1914 390
rect 1888 380 1890 382
rect 1894 381 1897 382
rect 1901 381 1904 382
rect 1894 380 1904 381
rect 1912 380 1914 382
rect 1922 389 1924 391
rect 1932 390 1942 391
rect 1932 389 1935 390
rect 1939 389 1942 390
rect 1946 389 1948 391
rect 1965 390 1969 398
rect 1922 381 1924 383
rect 1932 381 1942 383
rect 1946 381 1948 383
rect 1956 388 1958 390
rect 1962 388 1972 390
rect 1980 388 1982 390
rect 1897 365 1901 373
rect 1935 373 1939 381
rect 1956 380 1958 382
rect 1962 381 1965 382
rect 1969 381 1972 382
rect 1962 380 1972 381
rect 1980 380 1982 382
rect 1888 363 1890 365
rect 1894 363 1904 365
rect 1912 363 1914 365
rect 1888 355 1890 357
rect 1894 356 1897 357
rect 1901 356 1904 357
rect 1894 355 1904 356
rect 1912 355 1914 357
rect 1922 364 1924 366
rect 1932 365 1942 366
rect 1932 364 1935 365
rect 1939 364 1942 365
rect 1946 364 1948 366
rect 1965 365 1969 373
rect 1922 356 1924 358
rect 1932 356 1942 358
rect 1946 356 1948 358
rect 1956 363 1958 365
rect 1962 363 1972 365
rect 1980 363 1982 365
rect 1897 340 1901 348
rect 1935 348 1939 356
rect 1956 355 1958 357
rect 1962 356 1965 357
rect 1969 356 1972 357
rect 1962 355 1972 356
rect 1980 355 1982 357
rect 1888 338 1890 340
rect 1894 338 1904 340
rect 1912 338 1914 340
rect 1888 330 1890 332
rect 1894 331 1897 332
rect 1901 331 1904 332
rect 1894 330 1904 331
rect 1912 330 1914 332
rect 1922 339 1924 341
rect 1932 340 1942 341
rect 1932 339 1935 340
rect 1939 339 1942 340
rect 1946 339 1948 341
rect 1965 340 1969 348
rect 1922 331 1924 333
rect 1932 331 1942 333
rect 1946 331 1948 333
rect 1956 338 1958 340
rect 1962 338 1972 340
rect 1980 338 1982 340
rect 1897 315 1901 323
rect 1935 323 1939 331
rect 1956 330 1958 332
rect 1962 331 1965 332
rect 1969 331 1972 332
rect 1962 330 1972 331
rect 1980 330 1982 332
rect 1888 313 1890 315
rect 1894 313 1904 315
rect 1912 313 1914 315
rect 1888 305 1890 307
rect 1894 306 1897 307
rect 1901 306 1904 307
rect 1894 305 1904 306
rect 1912 305 1914 307
rect 1922 314 1924 316
rect 1932 315 1942 316
rect 1932 314 1935 315
rect 1939 314 1942 315
rect 1946 314 1948 316
rect 1965 315 1969 323
rect 1922 306 1924 308
rect 1932 306 1942 308
rect 1946 306 1948 308
rect 1956 313 1958 315
rect 1962 313 1972 315
rect 1980 313 1982 315
rect 1897 290 1901 298
rect 1935 298 1939 306
rect 1956 305 1958 307
rect 1962 306 1965 307
rect 1969 306 1972 307
rect 1962 305 1972 306
rect 1980 305 1982 307
rect 1888 288 1890 290
rect 1894 288 1904 290
rect 1912 288 1914 290
rect 1888 280 1890 282
rect 1894 281 1897 282
rect 1901 281 1904 282
rect 1894 280 1904 281
rect 1912 280 1914 282
rect 1922 289 1924 291
rect 1932 290 1942 291
rect 1932 289 1935 290
rect 1939 289 1942 290
rect 1946 289 1948 291
rect 1965 290 1969 298
rect 1922 281 1924 283
rect 1932 281 1942 283
rect 1946 281 1948 283
rect 1956 288 1958 290
rect 1962 288 1972 290
rect 1980 288 1982 290
rect 1897 265 1901 273
rect 1935 273 1939 281
rect 1956 280 1958 282
rect 1962 281 1965 282
rect 1969 281 1972 282
rect 1962 280 1972 281
rect 1980 280 1982 282
rect 1888 263 1890 265
rect 1894 263 1904 265
rect 1912 263 1914 265
rect 1888 255 1890 257
rect 1894 256 1897 257
rect 1901 256 1904 257
rect 1894 255 1904 256
rect 1912 255 1914 257
rect 1922 264 1924 266
rect 1932 265 1942 266
rect 1932 264 1935 265
rect 1939 264 1942 265
rect 1946 264 1948 266
rect 1965 265 1969 273
rect 1922 256 1924 258
rect 1932 256 1942 258
rect 1946 256 1948 258
rect 1956 263 1958 265
rect 1962 263 1972 265
rect 1980 263 1982 265
rect 1897 240 1901 248
rect 1935 248 1939 256
rect 1956 255 1958 257
rect 1962 256 1965 257
rect 1969 256 1972 257
rect 1962 255 1972 256
rect 1980 255 1982 257
rect 1888 238 1890 240
rect 1894 238 1904 240
rect 1912 238 1914 240
rect 1888 230 1890 232
rect 1894 231 1897 232
rect 1901 231 1904 232
rect 1894 230 1904 231
rect 1912 230 1914 232
rect 1922 239 1924 241
rect 1932 240 1942 241
rect 1932 239 1935 240
rect 1939 239 1942 240
rect 1946 239 1948 241
rect 1965 240 1969 248
rect 1922 231 1924 233
rect 1932 231 1942 233
rect 1946 231 1948 233
rect 1956 238 1958 240
rect 1962 238 1972 240
rect 1980 238 1982 240
rect 1897 215 1901 223
rect 1935 223 1939 231
rect 1956 230 1958 232
rect 1962 231 1965 232
rect 1969 231 1972 232
rect 1962 230 1972 231
rect 1980 230 1982 232
rect 1888 213 1890 215
rect 1894 213 1904 215
rect 1912 213 1914 215
rect 1888 205 1890 207
rect 1894 206 1897 207
rect 1901 206 1904 207
rect 1894 205 1904 206
rect 1912 205 1914 207
rect 1922 214 1924 216
rect 1932 215 1942 216
rect 1932 214 1935 215
rect 1939 214 1942 215
rect 1946 214 1948 216
rect 1965 215 1969 223
rect 1922 206 1924 208
rect 1932 206 1942 208
rect 1946 206 1948 208
rect 1956 213 1958 215
rect 1962 213 1972 215
rect 1980 213 1982 215
rect 1897 190 1901 198
rect 1935 198 1939 206
rect 1956 205 1958 207
rect 1962 206 1965 207
rect 1969 206 1972 207
rect 1962 205 1972 206
rect 1980 205 1982 207
rect 1888 188 1890 190
rect 1894 188 1904 190
rect 1912 188 1914 190
rect 1888 180 1890 182
rect 1894 181 1897 182
rect 1901 181 1904 182
rect 1894 180 1904 181
rect 1912 180 1914 182
rect 1922 189 1924 191
rect 1932 190 1942 191
rect 1932 189 1935 190
rect 1939 189 1942 190
rect 1946 189 1948 191
rect 1965 190 1969 198
rect 1922 181 1924 183
rect 1932 181 1942 183
rect 1946 181 1948 183
rect 1956 188 1958 190
rect 1962 188 1972 190
rect 1980 188 1982 190
rect 1897 165 1901 173
rect 1935 173 1939 181
rect 1956 180 1958 182
rect 1962 181 1965 182
rect 1969 181 1972 182
rect 1962 180 1972 181
rect 1980 180 1982 182
rect 1888 163 1890 165
rect 1894 163 1904 165
rect 1912 163 1914 165
rect 1888 155 1890 157
rect 1894 156 1897 157
rect 1901 156 1904 157
rect 1894 155 1904 156
rect 1912 155 1914 157
rect 1922 164 1924 166
rect 1932 165 1942 166
rect 1932 164 1935 165
rect 1939 164 1942 165
rect 1946 164 1948 166
rect 1965 165 1969 173
rect 1922 156 1924 158
rect 1932 156 1942 158
rect 1946 156 1948 158
rect 1956 163 1958 165
rect 1962 163 1972 165
rect 1980 163 1982 165
rect 1897 140 1901 148
rect 1935 148 1939 156
rect 1956 155 1958 157
rect 1962 156 1965 157
rect 1969 156 1972 157
rect 1962 155 1972 156
rect 1980 155 1982 157
rect 1888 138 1890 140
rect 1894 138 1904 140
rect 1912 138 1914 140
rect 1888 130 1890 132
rect 1894 131 1897 132
rect 1901 131 1904 132
rect 1894 130 1904 131
rect 1912 130 1914 132
rect 1922 139 1924 141
rect 1932 140 1942 141
rect 1932 139 1935 140
rect 1939 139 1942 140
rect 1946 139 1948 141
rect 1965 140 1969 148
rect 1922 131 1924 133
rect 1932 131 1942 133
rect 1946 131 1948 133
rect 1956 138 1958 140
rect 1962 138 1972 140
rect 1980 138 1982 140
rect 1897 115 1901 123
rect 1935 123 1939 131
rect 1956 130 1958 132
rect 1962 131 1965 132
rect 1969 131 1972 132
rect 1962 130 1972 131
rect 1980 130 1982 132
rect 1888 113 1890 115
rect 1894 113 1904 115
rect 1912 113 1914 115
rect 1888 105 1890 107
rect 1894 106 1897 107
rect 1901 106 1904 107
rect 1894 105 1904 106
rect 1912 105 1914 107
rect 1922 114 1924 116
rect 1932 115 1942 116
rect 1932 114 1935 115
rect 1939 114 1942 115
rect 1946 114 1948 116
rect 1965 115 1969 123
rect 1922 106 1924 108
rect 1932 106 1942 108
rect 1946 106 1948 108
rect 1956 113 1958 115
rect 1962 113 1972 115
rect 1980 113 1982 115
rect 1897 90 1901 98
rect 1935 98 1939 106
rect 1956 105 1958 107
rect 1962 106 1965 107
rect 1969 106 1972 107
rect 1962 105 1972 106
rect 1980 105 1982 107
rect 1888 88 1890 90
rect 1894 88 1904 90
rect 1912 88 1914 90
rect 1888 80 1890 82
rect 1894 81 1897 82
rect 1901 81 1904 82
rect 1894 80 1904 81
rect 1912 80 1914 82
rect 1922 89 1924 91
rect 1932 90 1942 91
rect 1932 89 1935 90
rect 1939 89 1942 90
rect 1946 89 1948 91
rect 1965 90 1969 98
rect 1922 81 1924 83
rect 1932 81 1942 83
rect 1946 81 1948 83
rect 1956 88 1958 90
rect 1962 88 1972 90
rect 1980 88 1982 90
rect 1897 65 1901 73
rect 1935 73 1939 81
rect 1956 80 1958 82
rect 1962 81 1965 82
rect 1969 81 1972 82
rect 1962 80 1972 81
rect 1980 80 1982 82
rect 1888 63 1890 65
rect 1894 63 1904 65
rect 1912 63 1914 65
rect 1888 55 1890 57
rect 1894 56 1897 57
rect 1901 56 1904 57
rect 1894 55 1904 56
rect 1912 55 1914 57
rect 1922 64 1924 66
rect 1932 65 1942 66
rect 1932 64 1935 65
rect 1939 64 1942 65
rect 1946 64 1948 66
rect 1965 65 1969 73
rect 1922 56 1924 58
rect 1932 56 1942 58
rect 1946 56 1948 58
rect 1956 63 1958 65
rect 1962 63 1972 65
rect 1980 63 1982 65
rect 1897 40 1901 48
rect 1935 48 1939 56
rect 1956 55 1958 57
rect 1962 56 1965 57
rect 1969 56 1972 57
rect 1962 55 1972 56
rect 1980 55 1982 57
rect 1888 38 1890 40
rect 1894 38 1904 40
rect 1912 38 1914 40
rect 1888 30 1890 32
rect 1894 31 1897 32
rect 1901 31 1904 32
rect 1894 30 1904 31
rect 1912 30 1914 32
rect 1922 39 1924 41
rect 1932 40 1942 41
rect 1932 39 1935 40
rect 1939 39 1942 40
rect 1946 39 1948 41
rect 1965 40 1969 48
rect 1922 31 1924 33
rect 1932 31 1942 33
rect 1946 31 1948 33
rect 1956 38 1958 40
rect 1962 38 1972 40
rect 1980 38 1982 40
rect 1935 23 1939 31
rect 1956 30 1958 32
rect 1962 31 1965 32
rect 1969 31 1972 32
rect 1962 30 1972 31
rect 1980 30 1982 32
rect 1897 21 1939 23
rect 1802 16 1807 17
rect 1966 16 1968 23
rect 1802 11 1968 16
<< ndiffusion >>
rect 1890 2015 1894 2016
rect 1942 2016 1946 2017
rect 1890 2012 1894 2013
rect 1890 2007 1894 2008
rect 1958 2015 1962 2016
rect 1942 2013 1946 2014
rect 1942 2008 1946 2009
rect 1958 2012 1962 2013
rect 1958 2007 1962 2008
rect 1890 2004 1894 2005
rect 1890 1990 1894 1991
rect 1942 2005 1946 2006
rect 1958 2004 1962 2005
rect 1942 1991 1946 1992
rect 1890 1987 1894 1988
rect 1890 1982 1894 1983
rect 1958 1990 1962 1991
rect 1942 1988 1946 1989
rect 1942 1983 1946 1984
rect 1958 1987 1962 1988
rect 1958 1982 1962 1983
rect 1890 1979 1894 1980
rect 1890 1965 1894 1966
rect 1942 1980 1946 1981
rect 1958 1979 1962 1980
rect 1942 1966 1946 1967
rect 1890 1962 1894 1963
rect 1890 1957 1894 1958
rect 1958 1965 1962 1966
rect 1942 1963 1946 1964
rect 1942 1958 1946 1959
rect 1958 1962 1962 1963
rect 1958 1957 1962 1958
rect 1890 1954 1894 1955
rect 1890 1940 1894 1941
rect 1942 1955 1946 1956
rect 1958 1954 1962 1955
rect 1942 1941 1946 1942
rect 1890 1937 1894 1938
rect 1890 1932 1894 1933
rect 1958 1940 1962 1941
rect 1942 1938 1946 1939
rect 1942 1933 1946 1934
rect 1958 1937 1962 1938
rect 1958 1932 1962 1933
rect 1890 1929 1894 1930
rect 1890 1915 1894 1916
rect 1942 1930 1946 1931
rect 1958 1929 1962 1930
rect 1942 1916 1946 1917
rect 1890 1912 1894 1913
rect 1890 1907 1894 1908
rect 1958 1915 1962 1916
rect 1942 1913 1946 1914
rect 1942 1908 1946 1909
rect 1958 1912 1962 1913
rect 1958 1907 1962 1908
rect 1890 1904 1894 1905
rect 1890 1890 1894 1891
rect 1942 1905 1946 1906
rect 1958 1904 1962 1905
rect 1942 1891 1946 1892
rect 1890 1887 1894 1888
rect 1890 1882 1894 1883
rect 1958 1890 1962 1891
rect 1942 1888 1946 1889
rect 1942 1883 1946 1884
rect 1958 1887 1962 1888
rect 1958 1882 1962 1883
rect 1890 1879 1894 1880
rect 1890 1865 1894 1866
rect 1942 1880 1946 1881
rect 1958 1879 1962 1880
rect 1942 1866 1946 1867
rect 1890 1862 1894 1863
rect 1890 1857 1894 1858
rect 1958 1865 1962 1866
rect 1942 1863 1946 1864
rect 1942 1858 1946 1859
rect 1958 1862 1962 1863
rect 1958 1857 1962 1858
rect 1890 1854 1894 1855
rect 1890 1840 1894 1841
rect 1942 1855 1946 1856
rect 1958 1854 1962 1855
rect 1942 1841 1946 1842
rect 1890 1837 1894 1838
rect 1890 1832 1894 1833
rect 1958 1840 1962 1841
rect 1942 1838 1946 1839
rect 1942 1833 1946 1834
rect 1958 1837 1962 1838
rect 1958 1832 1962 1833
rect 1890 1829 1894 1830
rect 1890 1815 1894 1816
rect 1942 1830 1946 1831
rect 1958 1829 1962 1830
rect 1942 1816 1946 1817
rect 1890 1812 1894 1813
rect 1890 1807 1894 1808
rect 1958 1815 1962 1816
rect 1942 1813 1946 1814
rect 1942 1808 1946 1809
rect 1958 1812 1962 1813
rect 1958 1807 1962 1808
rect 1890 1804 1894 1805
rect 1890 1790 1894 1791
rect 1942 1805 1946 1806
rect 1958 1804 1962 1805
rect 1942 1791 1946 1792
rect 1890 1787 1894 1788
rect 1890 1782 1894 1783
rect 1958 1790 1962 1791
rect 1942 1788 1946 1789
rect 1942 1783 1946 1784
rect 1958 1787 1962 1788
rect 1958 1782 1962 1783
rect 1890 1779 1894 1780
rect 1890 1765 1894 1766
rect 1942 1780 1946 1781
rect 1958 1779 1962 1780
rect 1942 1766 1946 1767
rect 1890 1762 1894 1763
rect 1890 1757 1894 1758
rect 1958 1765 1962 1766
rect 1942 1763 1946 1764
rect 1942 1758 1946 1759
rect 1958 1762 1962 1763
rect 1958 1757 1962 1758
rect 1890 1754 1894 1755
rect 1890 1740 1894 1741
rect 1942 1755 1946 1756
rect 1958 1754 1962 1755
rect 1942 1741 1946 1742
rect 1890 1737 1894 1738
rect 1890 1732 1894 1733
rect 1958 1740 1962 1741
rect 1942 1738 1946 1739
rect 1942 1733 1946 1734
rect 1958 1737 1962 1738
rect 1958 1732 1962 1733
rect 1890 1729 1894 1730
rect 1890 1715 1894 1716
rect 1942 1730 1946 1731
rect 1958 1729 1962 1730
rect 1942 1716 1946 1717
rect 1890 1712 1894 1713
rect 1890 1707 1894 1708
rect 1958 1715 1962 1716
rect 1942 1713 1946 1714
rect 1942 1708 1946 1709
rect 1958 1712 1962 1713
rect 1958 1707 1962 1708
rect 1890 1704 1894 1705
rect 1890 1690 1894 1691
rect 1942 1705 1946 1706
rect 1958 1704 1962 1705
rect 1942 1691 1946 1692
rect 1890 1687 1894 1688
rect 1890 1682 1894 1683
rect 1958 1690 1962 1691
rect 1942 1688 1946 1689
rect 1942 1683 1946 1684
rect 1958 1687 1962 1688
rect 1958 1682 1962 1683
rect 1890 1679 1894 1680
rect 1890 1665 1894 1666
rect 1942 1680 1946 1681
rect 1958 1679 1962 1680
rect 1942 1666 1946 1667
rect 1890 1662 1894 1663
rect 1890 1657 1894 1658
rect 1958 1665 1962 1666
rect 1942 1663 1946 1664
rect 1942 1658 1946 1659
rect 1958 1662 1962 1663
rect 1958 1657 1962 1658
rect 1890 1654 1894 1655
rect 1890 1640 1894 1641
rect 1942 1655 1946 1656
rect 1958 1654 1962 1655
rect 1942 1641 1946 1642
rect 1890 1637 1894 1638
rect 1890 1632 1894 1633
rect 1958 1640 1962 1641
rect 1942 1638 1946 1639
rect 1942 1633 1946 1634
rect 1958 1637 1962 1638
rect 1958 1632 1962 1633
rect 1890 1629 1894 1630
rect 1890 1615 1894 1616
rect 1942 1630 1946 1631
rect 1958 1629 1962 1630
rect 1942 1616 1946 1617
rect 1890 1612 1894 1613
rect 1890 1607 1894 1608
rect 1958 1615 1962 1616
rect 1942 1613 1946 1614
rect 1942 1608 1946 1609
rect 1958 1612 1962 1613
rect 1958 1607 1962 1608
rect 1890 1604 1894 1605
rect 1890 1590 1894 1591
rect 1942 1605 1946 1606
rect 1958 1604 1962 1605
rect 1942 1591 1946 1592
rect 1890 1587 1894 1588
rect 1890 1582 1894 1583
rect 1958 1590 1962 1591
rect 1942 1588 1946 1589
rect 1942 1583 1946 1584
rect 1958 1587 1962 1588
rect 1958 1582 1962 1583
rect 1890 1579 1894 1580
rect 1890 1565 1894 1566
rect 1942 1580 1946 1581
rect 1958 1579 1962 1580
rect 1942 1566 1946 1567
rect 1890 1562 1894 1563
rect 1890 1557 1894 1558
rect 1958 1565 1962 1566
rect 1942 1563 1946 1564
rect 1942 1558 1946 1559
rect 1958 1562 1962 1563
rect 1958 1557 1962 1558
rect 1890 1554 1894 1555
rect 1890 1540 1894 1541
rect 1942 1555 1946 1556
rect 1958 1554 1962 1555
rect 1942 1541 1946 1542
rect 1890 1537 1894 1538
rect 1890 1532 1894 1533
rect 1958 1540 1962 1541
rect 1942 1538 1946 1539
rect 1942 1533 1946 1534
rect 1958 1537 1962 1538
rect 1958 1532 1962 1533
rect 1890 1529 1894 1530
rect 1890 1515 1894 1516
rect 1942 1530 1946 1531
rect 1958 1529 1962 1530
rect 1942 1516 1946 1517
rect 1890 1512 1894 1513
rect 1890 1507 1894 1508
rect 1958 1515 1962 1516
rect 1942 1513 1946 1514
rect 1942 1508 1946 1509
rect 1958 1512 1962 1513
rect 1958 1507 1962 1508
rect 1890 1504 1894 1505
rect 1890 1490 1894 1491
rect 1942 1505 1946 1506
rect 1958 1504 1962 1505
rect 1942 1491 1946 1492
rect 1890 1487 1894 1488
rect 1890 1482 1894 1483
rect 1958 1490 1962 1491
rect 1942 1488 1946 1489
rect 1942 1483 1946 1484
rect 1958 1487 1962 1488
rect 1958 1482 1962 1483
rect 1890 1479 1894 1480
rect 1890 1465 1894 1466
rect 1942 1480 1946 1481
rect 1958 1479 1962 1480
rect 1942 1466 1946 1467
rect 1890 1462 1894 1463
rect 1890 1457 1894 1458
rect 1958 1465 1962 1466
rect 1942 1463 1946 1464
rect 1942 1458 1946 1459
rect 1958 1462 1962 1463
rect 1958 1457 1962 1458
rect 1890 1454 1894 1455
rect 1890 1440 1894 1441
rect 1942 1455 1946 1456
rect 1958 1454 1962 1455
rect 1942 1441 1946 1442
rect 1890 1437 1894 1438
rect 1890 1432 1894 1433
rect 1958 1440 1962 1441
rect 1942 1438 1946 1439
rect 1942 1433 1946 1434
rect 1958 1437 1962 1438
rect 1958 1432 1962 1433
rect 1890 1429 1894 1430
rect 1890 1415 1894 1416
rect 1942 1430 1946 1431
rect 1958 1429 1962 1430
rect 1942 1416 1946 1417
rect 1890 1412 1894 1413
rect 1890 1407 1894 1408
rect 1958 1415 1962 1416
rect 1942 1413 1946 1414
rect 1942 1408 1946 1409
rect 1958 1412 1962 1413
rect 1958 1407 1962 1408
rect 1890 1404 1894 1405
rect 1890 1390 1894 1391
rect 1942 1405 1946 1406
rect 1958 1404 1962 1405
rect 1942 1391 1946 1392
rect 1890 1387 1894 1388
rect 1890 1382 1894 1383
rect 1958 1390 1962 1391
rect 1942 1388 1946 1389
rect 1942 1383 1946 1384
rect 1958 1387 1962 1388
rect 1958 1382 1962 1383
rect 1756 1370 1758 1380
rect 1760 1370 1762 1380
rect 1890 1379 1894 1380
rect 1890 1365 1894 1366
rect 1942 1380 1946 1381
rect 1958 1379 1962 1380
rect 1942 1366 1946 1367
rect 1890 1362 1894 1363
rect 1890 1357 1894 1358
rect 1958 1365 1962 1366
rect 1942 1363 1946 1364
rect 1942 1358 1946 1359
rect 1958 1362 1962 1363
rect 1958 1357 1962 1358
rect 1890 1354 1894 1355
rect 1890 1340 1894 1341
rect 1942 1355 1946 1356
rect 1958 1354 1962 1355
rect 1942 1341 1946 1342
rect 1890 1337 1894 1338
rect 1890 1332 1894 1333
rect 1958 1340 1962 1341
rect 1942 1338 1946 1339
rect 1942 1333 1946 1334
rect 1958 1337 1962 1338
rect 1958 1332 1962 1333
rect 1890 1329 1894 1330
rect 1890 1315 1894 1316
rect 1942 1330 1946 1331
rect 1958 1329 1962 1330
rect 1942 1316 1946 1317
rect 1890 1312 1894 1313
rect 1890 1307 1894 1308
rect 1958 1315 1962 1316
rect 1942 1313 1946 1314
rect 1942 1308 1946 1309
rect 1958 1312 1962 1313
rect 1958 1307 1962 1308
rect 1890 1304 1894 1305
rect 1890 1290 1894 1291
rect 1942 1305 1946 1306
rect 1958 1304 1962 1305
rect 1942 1291 1946 1292
rect 1890 1287 1894 1288
rect 1890 1282 1894 1283
rect 1958 1290 1962 1291
rect 1942 1288 1946 1289
rect 1942 1283 1946 1284
rect 1958 1287 1962 1288
rect 1958 1282 1962 1283
rect 1890 1279 1894 1280
rect 1890 1265 1894 1266
rect 1942 1280 1946 1281
rect 1958 1279 1962 1280
rect 1942 1266 1946 1267
rect 1890 1262 1894 1263
rect 1890 1257 1894 1258
rect 1958 1265 1962 1266
rect 1942 1263 1946 1264
rect 1942 1258 1946 1259
rect 1958 1262 1962 1263
rect 1958 1257 1962 1258
rect 1890 1254 1894 1255
rect 1890 1240 1894 1241
rect 1942 1255 1946 1256
rect 1958 1254 1962 1255
rect 1942 1241 1946 1242
rect 1890 1237 1894 1238
rect 1890 1232 1894 1233
rect 1958 1240 1962 1241
rect 1942 1238 1946 1239
rect 1942 1233 1946 1234
rect 1958 1237 1962 1238
rect 1958 1232 1962 1233
rect 1890 1229 1894 1230
rect 1890 1215 1894 1216
rect 1942 1230 1946 1231
rect 1958 1229 1962 1230
rect 1942 1216 1946 1217
rect 1890 1212 1894 1213
rect 1890 1207 1894 1208
rect 1958 1215 1962 1216
rect 1942 1213 1946 1214
rect 1942 1208 1946 1209
rect 1958 1212 1962 1213
rect 1958 1207 1962 1208
rect 1890 1204 1894 1205
rect 910 1188 912 1198
rect 914 1188 916 1198
rect 1890 1190 1894 1191
rect 1942 1205 1946 1206
rect 1958 1204 1962 1205
rect 1942 1191 1946 1192
rect 1890 1187 1894 1188
rect 1890 1182 1894 1183
rect 1958 1190 1962 1191
rect 1942 1188 1946 1189
rect 1942 1183 1946 1184
rect 1958 1187 1962 1188
rect 1958 1182 1962 1183
rect 1890 1179 1894 1180
rect 1890 1165 1894 1166
rect 1942 1180 1946 1181
rect 1958 1179 1962 1180
rect 1942 1166 1946 1167
rect 1890 1162 1894 1163
rect 1890 1157 1894 1158
rect 1958 1165 1962 1166
rect 1942 1163 1946 1164
rect 1942 1158 1946 1159
rect 1958 1162 1962 1163
rect 1958 1157 1962 1158
rect 1890 1154 1894 1155
rect 1890 1140 1894 1141
rect 1942 1155 1946 1156
rect 1958 1154 1962 1155
rect 1942 1141 1946 1142
rect 1890 1137 1894 1138
rect 1890 1132 1894 1133
rect 1958 1140 1962 1141
rect 1942 1138 1946 1139
rect 1942 1133 1946 1134
rect 1958 1137 1962 1138
rect 1958 1132 1962 1133
rect 1890 1129 1894 1130
rect 1890 1115 1894 1116
rect 1942 1130 1946 1131
rect 1958 1129 1962 1130
rect 1942 1116 1946 1117
rect 1890 1112 1894 1113
rect 1890 1107 1894 1108
rect 1958 1115 1962 1116
rect 1942 1113 1946 1114
rect 1942 1108 1946 1109
rect 1958 1112 1962 1113
rect 1958 1107 1962 1108
rect 1890 1104 1894 1105
rect 1890 1090 1894 1091
rect 1942 1105 1946 1106
rect 1958 1104 1962 1105
rect 1942 1091 1946 1092
rect 1890 1087 1894 1088
rect 1890 1082 1894 1083
rect 1958 1090 1962 1091
rect 1942 1088 1946 1089
rect 1942 1083 1946 1084
rect 1958 1087 1962 1088
rect 1958 1082 1962 1083
rect 1890 1079 1894 1080
rect 1890 1065 1894 1066
rect 1942 1080 1946 1081
rect 1958 1079 1962 1080
rect 1942 1066 1946 1067
rect 1733 1055 1735 1065
rect 1737 1055 1739 1065
rect 1751 1055 1753 1065
rect 1755 1055 1757 1065
rect 1761 1055 1763 1065
rect 1765 1055 1767 1065
rect 1890 1062 1894 1063
rect 1890 1057 1894 1058
rect 1958 1065 1962 1066
rect 1942 1063 1946 1064
rect 1942 1058 1946 1059
rect 1958 1062 1962 1063
rect 1958 1057 1962 1058
rect 1890 1054 1894 1055
rect 1890 1040 1894 1041
rect 1942 1055 1946 1056
rect 1958 1054 1962 1055
rect 1942 1041 1946 1042
rect 1890 1037 1894 1038
rect 1890 1032 1894 1033
rect 1958 1040 1962 1041
rect 1942 1038 1946 1039
rect 1942 1033 1946 1034
rect 1958 1037 1962 1038
rect 1958 1032 1962 1033
rect 1890 1029 1894 1030
rect 1890 1015 1894 1016
rect 1942 1030 1946 1031
rect 1958 1029 1962 1030
rect 1942 1016 1946 1017
rect 1890 1012 1894 1013
rect 1890 1007 1894 1008
rect 1958 1015 1962 1016
rect 1942 1013 1946 1014
rect 1942 1008 1946 1009
rect 1958 1012 1962 1013
rect 1958 1007 1962 1008
rect 1890 1004 1894 1005
rect 1890 990 1894 991
rect 1942 1005 1946 1006
rect 1958 1004 1962 1005
rect 1942 991 1946 992
rect 1890 987 1894 988
rect 1890 982 1894 983
rect 1958 990 1962 991
rect 1942 988 1946 989
rect 1942 983 1946 984
rect 1958 987 1962 988
rect 1958 982 1962 983
rect 1890 979 1894 980
rect 1890 965 1894 966
rect 1942 980 1946 981
rect 1958 979 1962 980
rect 1942 966 1946 967
rect 1890 962 1894 963
rect 1890 957 1894 958
rect 1958 965 1962 966
rect 1942 963 1946 964
rect 1942 958 1946 959
rect 1958 962 1962 963
rect 1958 957 1962 958
rect 1890 954 1894 955
rect 1890 940 1894 941
rect 1942 955 1946 956
rect 1958 954 1962 955
rect 1942 941 1946 942
rect 1890 937 1894 938
rect 1890 932 1894 933
rect 1958 940 1962 941
rect 1942 938 1946 939
rect 1942 933 1946 934
rect 1958 937 1962 938
rect 1958 932 1962 933
rect 1890 929 1894 930
rect 1890 915 1894 916
rect 1942 930 1946 931
rect 1958 929 1962 930
rect 1942 916 1946 917
rect 1890 912 1894 913
rect 1890 907 1894 908
rect 1958 915 1962 916
rect 1942 913 1946 914
rect 1942 908 1946 909
rect 1958 912 1962 913
rect 1958 907 1962 908
rect 1890 904 1894 905
rect 1890 890 1894 891
rect 1942 905 1946 906
rect 1958 904 1962 905
rect 1942 891 1946 892
rect 1890 887 1894 888
rect 1890 882 1894 883
rect 1958 890 1962 891
rect 1942 888 1946 889
rect 1942 883 1946 884
rect 1958 887 1962 888
rect 1958 882 1962 883
rect 1890 879 1894 880
rect 1890 865 1894 866
rect 1942 880 1946 881
rect 1958 879 1962 880
rect 1942 866 1946 867
rect 1890 862 1894 863
rect 1890 857 1894 858
rect 1958 865 1962 866
rect 1942 863 1946 864
rect 1942 858 1946 859
rect 1958 862 1962 863
rect 1958 857 1962 858
rect 1890 854 1894 855
rect 1890 840 1894 841
rect 1942 855 1946 856
rect 1958 854 1962 855
rect 1942 841 1946 842
rect 1890 837 1894 838
rect 1890 832 1894 833
rect 1958 840 1962 841
rect 1942 838 1946 839
rect 1942 833 1946 834
rect 1958 837 1962 838
rect 1958 832 1962 833
rect 1890 829 1894 830
rect 1890 815 1894 816
rect 1942 830 1946 831
rect 1958 829 1962 830
rect 1942 816 1946 817
rect 1890 812 1894 813
rect 1890 807 1894 808
rect 1958 815 1962 816
rect 1942 813 1946 814
rect 1942 808 1946 809
rect 1958 812 1962 813
rect 1958 807 1962 808
rect 1890 804 1894 805
rect 1890 790 1894 791
rect 1942 805 1946 806
rect 1958 804 1962 805
rect 1942 791 1946 792
rect 1890 787 1894 788
rect 1890 782 1894 783
rect 1958 790 1962 791
rect 1942 788 1946 789
rect 1942 783 1946 784
rect 1958 787 1962 788
rect 1958 782 1962 783
rect 1890 779 1894 780
rect 1890 765 1894 766
rect 1942 780 1946 781
rect 1958 779 1962 780
rect 1942 766 1946 767
rect 1890 762 1894 763
rect 1890 757 1894 758
rect 1958 765 1962 766
rect 1942 763 1946 764
rect 1942 758 1946 759
rect 1958 762 1962 763
rect 1958 757 1962 758
rect 1890 754 1894 755
rect 1890 740 1894 741
rect 1942 755 1946 756
rect 1958 754 1962 755
rect 1942 741 1946 742
rect 1890 737 1894 738
rect 1890 732 1894 733
rect 1958 740 1962 741
rect 1942 738 1946 739
rect 1942 733 1946 734
rect 1958 737 1962 738
rect 1958 732 1962 733
rect 1890 729 1894 730
rect 1890 715 1894 716
rect 1942 730 1946 731
rect 1958 729 1962 730
rect 1942 716 1946 717
rect 1890 712 1894 713
rect 1890 707 1894 708
rect 1958 715 1962 716
rect 1942 713 1946 714
rect 1942 708 1946 709
rect 1958 712 1962 713
rect 1958 707 1962 708
rect 1890 704 1894 705
rect 1890 690 1894 691
rect 1942 705 1946 706
rect 1958 704 1962 705
rect 1942 691 1946 692
rect 1890 687 1894 688
rect 1890 682 1894 683
rect 1958 690 1962 691
rect 1942 688 1946 689
rect 1942 683 1946 684
rect 1958 687 1962 688
rect 1958 682 1962 683
rect 1890 679 1894 680
rect 1890 665 1894 666
rect 1942 680 1946 681
rect 1958 679 1962 680
rect 1942 666 1946 667
rect 1890 662 1894 663
rect 1890 657 1894 658
rect 1958 665 1962 666
rect 1942 663 1946 664
rect 1942 658 1946 659
rect 1958 662 1962 663
rect 1958 657 1962 658
rect 1890 654 1894 655
rect 1890 640 1894 641
rect 1942 655 1946 656
rect 1958 654 1962 655
rect 1942 641 1946 642
rect 1890 637 1894 638
rect 1890 632 1894 633
rect 1958 640 1962 641
rect 1942 638 1946 639
rect 1942 633 1946 634
rect 1958 637 1962 638
rect 1958 632 1962 633
rect 1890 629 1894 630
rect 1890 615 1894 616
rect 1942 630 1946 631
rect 1958 629 1962 630
rect 1942 616 1946 617
rect 1890 612 1894 613
rect 1890 607 1894 608
rect 1958 615 1962 616
rect 1942 613 1946 614
rect 1942 608 1946 609
rect 1958 612 1962 613
rect 1958 607 1962 608
rect 1890 604 1894 605
rect 1890 590 1894 591
rect 1942 605 1946 606
rect 1958 604 1962 605
rect 1942 591 1946 592
rect 1890 587 1894 588
rect 1890 582 1894 583
rect 1958 590 1962 591
rect 1942 588 1946 589
rect 1942 583 1946 584
rect 1958 587 1962 588
rect 1958 582 1962 583
rect 1890 579 1894 580
rect 1890 565 1894 566
rect 1942 580 1946 581
rect 1958 579 1962 580
rect 1942 566 1946 567
rect 1890 562 1894 563
rect 1890 557 1894 558
rect 1958 565 1962 566
rect 1942 563 1946 564
rect 1942 558 1946 559
rect 1958 562 1962 563
rect 1958 557 1962 558
rect 1890 554 1894 555
rect 1890 540 1894 541
rect 1942 555 1946 556
rect 1958 554 1962 555
rect 1942 541 1946 542
rect 1890 537 1894 538
rect 1890 532 1894 533
rect 1958 540 1962 541
rect 1942 538 1946 539
rect 1942 533 1946 534
rect 1958 537 1962 538
rect 1958 532 1962 533
rect 1890 529 1894 530
rect 1890 515 1894 516
rect 1942 530 1946 531
rect 1958 529 1962 530
rect 1942 516 1946 517
rect 1890 512 1894 513
rect 1890 507 1894 508
rect 1958 515 1962 516
rect 1942 513 1946 514
rect 1942 508 1946 509
rect 1958 512 1962 513
rect 1958 507 1962 508
rect 1890 504 1894 505
rect 1890 490 1894 491
rect 1942 505 1946 506
rect 1958 504 1962 505
rect 1942 491 1946 492
rect 1890 487 1894 488
rect 1890 482 1894 483
rect 1958 490 1962 491
rect 1942 488 1946 489
rect 1942 483 1946 484
rect 1958 487 1962 488
rect 1958 482 1962 483
rect 1890 479 1894 480
rect 1890 465 1894 466
rect 1942 480 1946 481
rect 1958 479 1962 480
rect 1942 466 1946 467
rect 1890 462 1894 463
rect 1890 457 1894 458
rect 1958 465 1962 466
rect 1942 463 1946 464
rect 1942 458 1946 459
rect 1958 462 1962 463
rect 1958 457 1962 458
rect 1890 454 1894 455
rect 1890 440 1894 441
rect 1942 455 1946 456
rect 1958 454 1962 455
rect 1942 441 1946 442
rect 1890 437 1894 438
rect 1890 432 1894 433
rect 1958 440 1962 441
rect 1942 438 1946 439
rect 1942 433 1946 434
rect 1958 437 1962 438
rect 1958 432 1962 433
rect 1890 429 1894 430
rect 1890 415 1894 416
rect 1942 430 1946 431
rect 1958 429 1962 430
rect 1942 416 1946 417
rect 1890 412 1894 413
rect 1890 407 1894 408
rect 1958 415 1962 416
rect 1942 413 1946 414
rect 1942 408 1946 409
rect 1958 412 1962 413
rect 1958 407 1962 408
rect 1890 404 1894 405
rect 1890 390 1894 391
rect 1942 405 1946 406
rect 1958 404 1962 405
rect 1942 391 1946 392
rect 1890 387 1894 388
rect 1890 382 1894 383
rect 1958 390 1962 391
rect 1942 388 1946 389
rect 1942 383 1946 384
rect 1958 387 1962 388
rect 1958 382 1962 383
rect 1890 379 1894 380
rect 1890 365 1894 366
rect 1942 380 1946 381
rect 1958 379 1962 380
rect 1942 366 1946 367
rect 1890 362 1894 363
rect 1890 357 1894 358
rect 1958 365 1962 366
rect 1942 363 1946 364
rect 1942 358 1946 359
rect 1958 362 1962 363
rect 1958 357 1962 358
rect 1890 354 1894 355
rect 1890 340 1894 341
rect 1942 355 1946 356
rect 1958 354 1962 355
rect 1942 341 1946 342
rect 1890 337 1894 338
rect 1890 332 1894 333
rect 1958 340 1962 341
rect 1942 338 1946 339
rect 1942 333 1946 334
rect 1958 337 1962 338
rect 1958 332 1962 333
rect 1890 329 1894 330
rect 1890 315 1894 316
rect 1942 330 1946 331
rect 1958 329 1962 330
rect 1942 316 1946 317
rect 1890 312 1894 313
rect 1890 307 1894 308
rect 1958 315 1962 316
rect 1942 313 1946 314
rect 1942 308 1946 309
rect 1958 312 1962 313
rect 1958 307 1962 308
rect 1890 304 1894 305
rect 1890 290 1894 291
rect 1942 305 1946 306
rect 1958 304 1962 305
rect 1942 291 1946 292
rect 1890 287 1894 288
rect 1890 282 1894 283
rect 1958 290 1962 291
rect 1942 288 1946 289
rect 1942 283 1946 284
rect 1958 287 1962 288
rect 1958 282 1962 283
rect 1890 279 1894 280
rect 1890 265 1894 266
rect 1942 280 1946 281
rect 1958 279 1962 280
rect 1942 266 1946 267
rect 1890 262 1894 263
rect 1890 257 1894 258
rect 1958 265 1962 266
rect 1942 263 1946 264
rect 1942 258 1946 259
rect 1958 262 1962 263
rect 1958 257 1962 258
rect 1890 254 1894 255
rect 1890 240 1894 241
rect 1942 255 1946 256
rect 1958 254 1962 255
rect 1942 241 1946 242
rect 1890 237 1894 238
rect 1890 232 1894 233
rect 1958 240 1962 241
rect 1942 238 1946 239
rect 1942 233 1946 234
rect 1958 237 1962 238
rect 1958 232 1962 233
rect 1890 229 1894 230
rect 1890 215 1894 216
rect 1942 230 1946 231
rect 1958 229 1962 230
rect 1942 216 1946 217
rect 1890 212 1894 213
rect 1890 207 1894 208
rect 1958 215 1962 216
rect 1942 213 1946 214
rect 1942 208 1946 209
rect 1958 212 1962 213
rect 1958 207 1962 208
rect 1890 204 1894 205
rect 1890 190 1894 191
rect 1942 205 1946 206
rect 1958 204 1962 205
rect 1942 191 1946 192
rect 1890 187 1894 188
rect 1890 182 1894 183
rect 1958 190 1962 191
rect 1942 188 1946 189
rect 1942 183 1946 184
rect 1958 187 1962 188
rect 1958 182 1962 183
rect 1890 179 1894 180
rect 1890 165 1894 166
rect 1942 180 1946 181
rect 1958 179 1962 180
rect 1942 166 1946 167
rect 1890 162 1894 163
rect 1890 157 1894 158
rect 1958 165 1962 166
rect 1942 163 1946 164
rect 1942 158 1946 159
rect 1958 162 1962 163
rect 1958 157 1962 158
rect 1890 154 1894 155
rect 1890 140 1894 141
rect 1942 155 1946 156
rect 1958 154 1962 155
rect 1942 141 1946 142
rect 1890 137 1894 138
rect 1890 132 1894 133
rect 1958 140 1962 141
rect 1942 138 1946 139
rect 1942 133 1946 134
rect 1958 137 1962 138
rect 1958 132 1962 133
rect 1890 129 1894 130
rect 1890 115 1894 116
rect 1942 130 1946 131
rect 1958 129 1962 130
rect 1942 116 1946 117
rect 1890 112 1894 113
rect 1890 107 1894 108
rect 1958 115 1962 116
rect 1942 113 1946 114
rect 1942 108 1946 109
rect 1958 112 1962 113
rect 1958 107 1962 108
rect 1890 104 1894 105
rect 1890 90 1894 91
rect 1942 105 1946 106
rect 1958 104 1962 105
rect 1942 91 1946 92
rect 1890 87 1894 88
rect 1890 82 1894 83
rect 1958 90 1962 91
rect 1942 88 1946 89
rect 1942 83 1946 84
rect 1958 87 1962 88
rect 1958 82 1962 83
rect 1890 79 1894 80
rect 1890 65 1894 66
rect 1942 80 1946 81
rect 1958 79 1962 80
rect 1942 66 1946 67
rect 1890 62 1894 63
rect 1890 57 1894 58
rect 1958 65 1962 66
rect 1942 63 1946 64
rect 1942 58 1946 59
rect 1958 62 1962 63
rect 1958 57 1962 58
rect 1890 54 1894 55
rect 1890 40 1894 41
rect 1942 55 1946 56
rect 1958 54 1962 55
rect 1942 41 1946 42
rect 1890 37 1894 38
rect 1890 32 1894 33
rect 1958 40 1962 41
rect 1942 38 1946 39
rect 1942 33 1946 34
rect 1958 37 1962 38
rect 1958 32 1962 33
rect 1890 29 1894 30
rect 1942 30 1946 31
rect 1958 29 1962 30
<< pdiffusion >>
rect 1924 2016 1932 2017
rect 1904 2015 1912 2016
rect 1904 2012 1912 2013
rect 1904 2007 1912 2008
rect 1924 2013 1932 2014
rect 1972 2015 1980 2016
rect 1924 2008 1932 2009
rect 1972 2012 1980 2013
rect 1924 2005 1932 2006
rect 1904 2004 1912 2005
rect 1972 2007 1980 2008
rect 1972 2004 1980 2005
rect 1924 1991 1932 1992
rect 1904 1990 1912 1991
rect 1904 1987 1912 1988
rect 1904 1982 1912 1983
rect 1924 1988 1932 1989
rect 1972 1990 1980 1991
rect 1924 1983 1932 1984
rect 1972 1987 1980 1988
rect 1924 1980 1932 1981
rect 1904 1979 1912 1980
rect 1972 1982 1980 1983
rect 1972 1979 1980 1980
rect 1924 1966 1932 1967
rect 1904 1965 1912 1966
rect 1904 1962 1912 1963
rect 1904 1957 1912 1958
rect 1924 1963 1932 1964
rect 1972 1965 1980 1966
rect 1924 1958 1932 1959
rect 1972 1962 1980 1963
rect 1924 1955 1932 1956
rect 1904 1954 1912 1955
rect 1972 1957 1980 1958
rect 1972 1954 1980 1955
rect 1924 1941 1932 1942
rect 1904 1940 1912 1941
rect 1904 1937 1912 1938
rect 1904 1932 1912 1933
rect 1924 1938 1932 1939
rect 1972 1940 1980 1941
rect 1924 1933 1932 1934
rect 1972 1937 1980 1938
rect 1924 1930 1932 1931
rect 1904 1929 1912 1930
rect 1972 1932 1980 1933
rect 1972 1929 1980 1930
rect 1924 1916 1932 1917
rect 1904 1915 1912 1916
rect 1904 1912 1912 1913
rect 1904 1907 1912 1908
rect 1924 1913 1932 1914
rect 1972 1915 1980 1916
rect 1924 1908 1932 1909
rect 1972 1912 1980 1913
rect 1924 1905 1932 1906
rect 1904 1904 1912 1905
rect 1972 1907 1980 1908
rect 1972 1904 1980 1905
rect 1924 1891 1932 1892
rect 1904 1890 1912 1891
rect 1904 1887 1912 1888
rect 1904 1882 1912 1883
rect 1924 1888 1932 1889
rect 1972 1890 1980 1891
rect 1924 1883 1932 1884
rect 1972 1887 1980 1888
rect 1924 1880 1932 1881
rect 1904 1879 1912 1880
rect 1972 1882 1980 1883
rect 1972 1879 1980 1880
rect 1924 1866 1932 1867
rect 1904 1865 1912 1866
rect 1904 1862 1912 1863
rect 1904 1857 1912 1858
rect 1924 1863 1932 1864
rect 1972 1865 1980 1866
rect 1924 1858 1932 1859
rect 1972 1862 1980 1863
rect 1924 1855 1932 1856
rect 1904 1854 1912 1855
rect 1972 1857 1980 1858
rect 1972 1854 1980 1855
rect 1924 1841 1932 1842
rect 1904 1840 1912 1841
rect 1904 1837 1912 1838
rect 1904 1832 1912 1833
rect 1924 1838 1932 1839
rect 1972 1840 1980 1841
rect 1924 1833 1932 1834
rect 1972 1837 1980 1838
rect 1924 1830 1932 1831
rect 1904 1829 1912 1830
rect 1972 1832 1980 1833
rect 1972 1829 1980 1830
rect 1924 1816 1932 1817
rect 1904 1815 1912 1816
rect 1904 1812 1912 1813
rect 1904 1807 1912 1808
rect 1924 1813 1932 1814
rect 1972 1815 1980 1816
rect 1924 1808 1932 1809
rect 1972 1812 1980 1813
rect 1924 1805 1932 1806
rect 1904 1804 1912 1805
rect 1972 1807 1980 1808
rect 1972 1804 1980 1805
rect 1924 1791 1932 1792
rect 1904 1790 1912 1791
rect 1904 1787 1912 1788
rect 1904 1782 1912 1783
rect 1924 1788 1932 1789
rect 1972 1790 1980 1791
rect 1924 1783 1932 1784
rect 1972 1787 1980 1788
rect 1924 1780 1932 1781
rect 1904 1779 1912 1780
rect 1972 1782 1980 1783
rect 1972 1779 1980 1780
rect 1924 1766 1932 1767
rect 1904 1765 1912 1766
rect 1904 1762 1912 1763
rect 1904 1757 1912 1758
rect 1924 1763 1932 1764
rect 1972 1765 1980 1766
rect 1924 1758 1932 1759
rect 1972 1762 1980 1763
rect 1924 1755 1932 1756
rect 1904 1754 1912 1755
rect 1972 1757 1980 1758
rect 1972 1754 1980 1755
rect 1924 1741 1932 1742
rect 1904 1740 1912 1741
rect 1904 1737 1912 1738
rect 1904 1732 1912 1733
rect 1924 1738 1932 1739
rect 1972 1740 1980 1741
rect 1924 1733 1932 1734
rect 1972 1737 1980 1738
rect 1924 1730 1932 1731
rect 1904 1729 1912 1730
rect 1972 1732 1980 1733
rect 1972 1729 1980 1730
rect 1924 1716 1932 1717
rect 1904 1715 1912 1716
rect 1904 1712 1912 1713
rect 1904 1707 1912 1708
rect 1924 1713 1932 1714
rect 1972 1715 1980 1716
rect 1924 1708 1932 1709
rect 1972 1712 1980 1713
rect 1924 1705 1932 1706
rect 1904 1704 1912 1705
rect 1972 1707 1980 1708
rect 1972 1704 1980 1705
rect 1924 1691 1932 1692
rect 1904 1690 1912 1691
rect 1904 1687 1912 1688
rect 1904 1682 1912 1683
rect 1924 1688 1932 1689
rect 1972 1690 1980 1691
rect 1924 1683 1932 1684
rect 1972 1687 1980 1688
rect 1924 1680 1932 1681
rect 1904 1679 1912 1680
rect 1972 1682 1980 1683
rect 1972 1679 1980 1680
rect 1924 1666 1932 1667
rect 1904 1665 1912 1666
rect 1904 1662 1912 1663
rect 1904 1657 1912 1658
rect 1924 1663 1932 1664
rect 1972 1665 1980 1666
rect 1924 1658 1932 1659
rect 1972 1662 1980 1663
rect 1924 1655 1932 1656
rect 1904 1654 1912 1655
rect 1972 1657 1980 1658
rect 1972 1654 1980 1655
rect 1924 1641 1932 1642
rect 1904 1640 1912 1641
rect 1904 1637 1912 1638
rect 1904 1632 1912 1633
rect 1924 1638 1932 1639
rect 1972 1640 1980 1641
rect 1924 1633 1932 1634
rect 1972 1637 1980 1638
rect 1924 1630 1932 1631
rect 1904 1629 1912 1630
rect 1972 1632 1980 1633
rect 1972 1629 1980 1630
rect 1924 1616 1932 1617
rect 1904 1615 1912 1616
rect 1904 1612 1912 1613
rect 1904 1607 1912 1608
rect 1924 1613 1932 1614
rect 1972 1615 1980 1616
rect 1924 1608 1932 1609
rect 1972 1612 1980 1613
rect 1924 1605 1932 1606
rect 1904 1604 1912 1605
rect 1972 1607 1980 1608
rect 1972 1604 1980 1605
rect 1924 1591 1932 1592
rect 1904 1590 1912 1591
rect 1904 1587 1912 1588
rect 1904 1582 1912 1583
rect 1924 1588 1932 1589
rect 1972 1590 1980 1591
rect 1924 1583 1932 1584
rect 1972 1587 1980 1588
rect 1924 1580 1932 1581
rect 1904 1579 1912 1580
rect 1972 1582 1980 1583
rect 1972 1579 1980 1580
rect 1924 1566 1932 1567
rect 1904 1565 1912 1566
rect 1904 1562 1912 1563
rect 1904 1557 1912 1558
rect 1924 1563 1932 1564
rect 1972 1565 1980 1566
rect 1924 1558 1932 1559
rect 1972 1562 1980 1563
rect 1924 1555 1932 1556
rect 1904 1554 1912 1555
rect 1972 1557 1980 1558
rect 1972 1554 1980 1555
rect 1924 1541 1932 1542
rect 1904 1540 1912 1541
rect 1904 1537 1912 1538
rect 1904 1532 1912 1533
rect 1924 1538 1932 1539
rect 1972 1540 1980 1541
rect 1924 1533 1932 1534
rect 1972 1537 1980 1538
rect 1924 1530 1932 1531
rect 1904 1529 1912 1530
rect 1972 1532 1980 1533
rect 1972 1529 1980 1530
rect 1924 1516 1932 1517
rect 1904 1515 1912 1516
rect 1904 1512 1912 1513
rect 1904 1507 1912 1508
rect 1924 1513 1932 1514
rect 1972 1515 1980 1516
rect 1924 1508 1932 1509
rect 1972 1512 1980 1513
rect 1924 1505 1932 1506
rect 1904 1504 1912 1505
rect 1972 1507 1980 1508
rect 1972 1504 1980 1505
rect 1924 1491 1932 1492
rect 1904 1490 1912 1491
rect 1904 1487 1912 1488
rect 1904 1482 1912 1483
rect 1924 1488 1932 1489
rect 1972 1490 1980 1491
rect 1924 1483 1932 1484
rect 1972 1487 1980 1488
rect 1924 1480 1932 1481
rect 1904 1479 1912 1480
rect 1972 1482 1980 1483
rect 1972 1479 1980 1480
rect 1924 1466 1932 1467
rect 1904 1465 1912 1466
rect 1904 1462 1912 1463
rect 1904 1457 1912 1458
rect 1924 1463 1932 1464
rect 1972 1465 1980 1466
rect 1924 1458 1932 1459
rect 1972 1462 1980 1463
rect 1924 1455 1932 1456
rect 1904 1454 1912 1455
rect 1972 1457 1980 1458
rect 1972 1454 1980 1455
rect 1924 1441 1932 1442
rect 1904 1440 1912 1441
rect 1904 1437 1912 1438
rect 1904 1432 1912 1433
rect 1924 1438 1932 1439
rect 1972 1440 1980 1441
rect 1924 1433 1932 1434
rect 1972 1437 1980 1438
rect 1924 1430 1932 1431
rect 1904 1429 1912 1430
rect 1972 1432 1980 1433
rect 1972 1429 1980 1430
rect 1924 1416 1932 1417
rect 1904 1415 1912 1416
rect 1756 1390 1758 1410
rect 1760 1390 1762 1410
rect 1904 1412 1912 1413
rect 1904 1407 1912 1408
rect 1924 1413 1932 1414
rect 1972 1415 1980 1416
rect 1924 1408 1932 1409
rect 1972 1412 1980 1413
rect 1924 1405 1932 1406
rect 1904 1404 1912 1405
rect 1972 1407 1980 1408
rect 1972 1404 1980 1405
rect 1924 1391 1932 1392
rect 1904 1390 1912 1391
rect 1904 1387 1912 1388
rect 1904 1382 1912 1383
rect 1924 1388 1932 1389
rect 1972 1390 1980 1391
rect 1924 1383 1932 1384
rect 1972 1387 1980 1388
rect 1924 1380 1932 1381
rect 1904 1379 1912 1380
rect 1972 1382 1980 1383
rect 1972 1379 1980 1380
rect 1924 1366 1932 1367
rect 1904 1365 1912 1366
rect 1904 1362 1912 1363
rect 1904 1357 1912 1358
rect 1924 1363 1932 1364
rect 1972 1365 1980 1366
rect 1924 1358 1932 1359
rect 1972 1362 1980 1363
rect 1924 1355 1932 1356
rect 1904 1354 1912 1355
rect 1972 1357 1980 1358
rect 1972 1354 1980 1355
rect 1924 1341 1932 1342
rect 1904 1340 1912 1341
rect 1904 1337 1912 1338
rect 1904 1332 1912 1333
rect 1924 1338 1932 1339
rect 1972 1340 1980 1341
rect 1924 1333 1932 1334
rect 1972 1337 1980 1338
rect 1924 1330 1932 1331
rect 1904 1329 1912 1330
rect 1972 1332 1980 1333
rect 1972 1329 1980 1330
rect 1924 1316 1932 1317
rect 1904 1315 1912 1316
rect 1904 1312 1912 1313
rect 1904 1307 1912 1308
rect 1924 1313 1932 1314
rect 1972 1315 1980 1316
rect 1924 1308 1932 1309
rect 1972 1312 1980 1313
rect 1924 1305 1932 1306
rect 1904 1304 1912 1305
rect 1972 1307 1980 1308
rect 1972 1304 1980 1305
rect 1924 1291 1932 1292
rect 1904 1290 1912 1291
rect 1904 1287 1912 1288
rect 1904 1282 1912 1283
rect 1924 1288 1932 1289
rect 1972 1290 1980 1291
rect 1924 1283 1932 1284
rect 1972 1287 1980 1288
rect 1924 1280 1932 1281
rect 1904 1279 1912 1280
rect 1972 1282 1980 1283
rect 1972 1279 1980 1280
rect 1924 1266 1932 1267
rect 1904 1265 1912 1266
rect 1904 1262 1912 1263
rect 1904 1257 1912 1258
rect 1924 1263 1932 1264
rect 1972 1265 1980 1266
rect 1924 1258 1932 1259
rect 1972 1262 1980 1263
rect 1924 1255 1932 1256
rect 1904 1254 1912 1255
rect 1972 1257 1980 1258
rect 1972 1254 1980 1255
rect 1924 1241 1932 1242
rect 1904 1240 1912 1241
rect 1904 1237 1912 1238
rect 1904 1232 1912 1233
rect 1924 1238 1932 1239
rect 1972 1240 1980 1241
rect 1924 1233 1932 1234
rect 1972 1237 1980 1238
rect 1924 1230 1932 1231
rect 1904 1229 1912 1230
rect 1972 1232 1980 1233
rect 1972 1229 1980 1230
rect 1924 1216 1932 1217
rect 1904 1215 1912 1216
rect 1904 1212 1912 1213
rect 1904 1207 1912 1208
rect 1924 1213 1932 1214
rect 1972 1215 1980 1216
rect 1924 1208 1932 1209
rect 1972 1212 1980 1213
rect 1924 1205 1932 1206
rect 1904 1204 1912 1205
rect 1972 1207 1980 1208
rect 1972 1204 1980 1205
rect 1924 1191 1932 1192
rect 1904 1190 1912 1191
rect 1904 1187 1912 1188
rect 1904 1182 1912 1183
rect 1924 1188 1932 1189
rect 1972 1190 1980 1191
rect 1924 1183 1932 1184
rect 1972 1187 1980 1188
rect 1924 1180 1932 1181
rect 910 1158 912 1178
rect 914 1158 916 1178
rect 1904 1179 1912 1180
rect 1972 1182 1980 1183
rect 1972 1179 1980 1180
rect 1924 1166 1932 1167
rect 1904 1165 1912 1166
rect 1904 1162 1912 1163
rect 1904 1157 1912 1158
rect 1924 1163 1932 1164
rect 1972 1165 1980 1166
rect 1924 1158 1932 1159
rect 1972 1162 1980 1163
rect 1924 1155 1932 1156
rect 1904 1154 1912 1155
rect 1972 1157 1980 1158
rect 1972 1154 1980 1155
rect 1924 1141 1932 1142
rect 1904 1140 1912 1141
rect 1904 1137 1912 1138
rect 1904 1132 1912 1133
rect 1924 1138 1932 1139
rect 1972 1140 1980 1141
rect 1924 1133 1932 1134
rect 1972 1137 1980 1138
rect 1924 1130 1932 1131
rect 1904 1129 1912 1130
rect 1972 1132 1980 1133
rect 1972 1129 1980 1130
rect 1924 1116 1932 1117
rect 1904 1115 1912 1116
rect 1904 1112 1912 1113
rect 1904 1107 1912 1108
rect 1924 1113 1932 1114
rect 1972 1115 1980 1116
rect 1924 1108 1932 1109
rect 1972 1112 1980 1113
rect 1924 1105 1932 1106
rect 1904 1104 1912 1105
rect 1733 1075 1735 1093
rect 1737 1075 1739 1093
rect 1751 1075 1753 1093
rect 1755 1075 1757 1093
rect 1761 1075 1763 1093
rect 1765 1075 1767 1093
rect 1972 1107 1980 1108
rect 1972 1104 1980 1105
rect 1924 1091 1932 1092
rect 1904 1090 1912 1091
rect 1904 1087 1912 1088
rect 1904 1082 1912 1083
rect 1924 1088 1932 1089
rect 1972 1090 1980 1091
rect 1924 1083 1932 1084
rect 1972 1087 1980 1088
rect 1924 1080 1932 1081
rect 1904 1079 1912 1080
rect 1972 1082 1980 1083
rect 1972 1079 1980 1080
rect 1924 1066 1932 1067
rect 1904 1065 1912 1066
rect 1904 1062 1912 1063
rect 1904 1057 1912 1058
rect 1924 1063 1932 1064
rect 1972 1065 1980 1066
rect 1924 1058 1932 1059
rect 1972 1062 1980 1063
rect 1924 1055 1932 1056
rect 1904 1054 1912 1055
rect 1972 1057 1980 1058
rect 1972 1054 1980 1055
rect 1924 1041 1932 1042
rect 1904 1040 1912 1041
rect 1904 1037 1912 1038
rect 1904 1032 1912 1033
rect 1924 1038 1932 1039
rect 1972 1040 1980 1041
rect 1924 1033 1932 1034
rect 1972 1037 1980 1038
rect 1924 1030 1932 1031
rect 1904 1029 1912 1030
rect 1972 1032 1980 1033
rect 1972 1029 1980 1030
rect 1924 1016 1932 1017
rect 1904 1015 1912 1016
rect 1904 1012 1912 1013
rect 1904 1007 1912 1008
rect 1924 1013 1932 1014
rect 1972 1015 1980 1016
rect 1924 1008 1932 1009
rect 1972 1012 1980 1013
rect 1924 1005 1932 1006
rect 1904 1004 1912 1005
rect 1972 1007 1980 1008
rect 1972 1004 1980 1005
rect 1924 991 1932 992
rect 1904 990 1912 991
rect 1904 987 1912 988
rect 1904 982 1912 983
rect 1924 988 1932 989
rect 1972 990 1980 991
rect 1924 983 1932 984
rect 1972 987 1980 988
rect 1924 980 1932 981
rect 1904 979 1912 980
rect 1972 982 1980 983
rect 1972 979 1980 980
rect 1924 966 1932 967
rect 1904 965 1912 966
rect 1904 962 1912 963
rect 1904 957 1912 958
rect 1924 963 1932 964
rect 1972 965 1980 966
rect 1924 958 1932 959
rect 1972 962 1980 963
rect 1924 955 1932 956
rect 1904 954 1912 955
rect 1972 957 1980 958
rect 1972 954 1980 955
rect 1924 941 1932 942
rect 1904 940 1912 941
rect 1904 937 1912 938
rect 1904 932 1912 933
rect 1924 938 1932 939
rect 1972 940 1980 941
rect 1924 933 1932 934
rect 1972 937 1980 938
rect 1924 930 1932 931
rect 1904 929 1912 930
rect 1972 932 1980 933
rect 1972 929 1980 930
rect 1924 916 1932 917
rect 1904 915 1912 916
rect 1904 912 1912 913
rect 1904 907 1912 908
rect 1924 913 1932 914
rect 1972 915 1980 916
rect 1924 908 1932 909
rect 1972 912 1980 913
rect 1924 905 1932 906
rect 1904 904 1912 905
rect 1972 907 1980 908
rect 1972 904 1980 905
rect 1924 891 1932 892
rect 1904 890 1912 891
rect 1904 887 1912 888
rect 1904 882 1912 883
rect 1924 888 1932 889
rect 1972 890 1980 891
rect 1924 883 1932 884
rect 1972 887 1980 888
rect 1924 880 1932 881
rect 1904 879 1912 880
rect 1972 882 1980 883
rect 1972 879 1980 880
rect 1924 866 1932 867
rect 1904 865 1912 866
rect 1904 862 1912 863
rect 1904 857 1912 858
rect 1924 863 1932 864
rect 1972 865 1980 866
rect 1924 858 1932 859
rect 1972 862 1980 863
rect 1924 855 1932 856
rect 1904 854 1912 855
rect 1972 857 1980 858
rect 1972 854 1980 855
rect 1924 841 1932 842
rect 1904 840 1912 841
rect 1904 837 1912 838
rect 1904 832 1912 833
rect 1924 838 1932 839
rect 1972 840 1980 841
rect 1924 833 1932 834
rect 1972 837 1980 838
rect 1924 830 1932 831
rect 1904 829 1912 830
rect 1972 832 1980 833
rect 1972 829 1980 830
rect 1924 816 1932 817
rect 1904 815 1912 816
rect 1904 812 1912 813
rect 1904 807 1912 808
rect 1924 813 1932 814
rect 1972 815 1980 816
rect 1924 808 1932 809
rect 1972 812 1980 813
rect 1924 805 1932 806
rect 1904 804 1912 805
rect 1972 807 1980 808
rect 1972 804 1980 805
rect 1924 791 1932 792
rect 1904 790 1912 791
rect 1904 787 1912 788
rect 1904 782 1912 783
rect 1924 788 1932 789
rect 1972 790 1980 791
rect 1924 783 1932 784
rect 1972 787 1980 788
rect 1924 780 1932 781
rect 1904 779 1912 780
rect 1972 782 1980 783
rect 1972 779 1980 780
rect 1924 766 1932 767
rect 1904 765 1912 766
rect 1904 762 1912 763
rect 1904 757 1912 758
rect 1924 763 1932 764
rect 1972 765 1980 766
rect 1924 758 1932 759
rect 1972 762 1980 763
rect 1924 755 1932 756
rect 1904 754 1912 755
rect 1972 757 1980 758
rect 1972 754 1980 755
rect 1924 741 1932 742
rect 1904 740 1912 741
rect 1904 737 1912 738
rect 1904 732 1912 733
rect 1924 738 1932 739
rect 1972 740 1980 741
rect 1924 733 1932 734
rect 1972 737 1980 738
rect 1924 730 1932 731
rect 1904 729 1912 730
rect 1972 732 1980 733
rect 1972 729 1980 730
rect 1924 716 1932 717
rect 1904 715 1912 716
rect 1904 712 1912 713
rect 1904 707 1912 708
rect 1924 713 1932 714
rect 1972 715 1980 716
rect 1924 708 1932 709
rect 1972 712 1980 713
rect 1924 705 1932 706
rect 1904 704 1912 705
rect 1972 707 1980 708
rect 1972 704 1980 705
rect 1924 691 1932 692
rect 1904 690 1912 691
rect 1904 687 1912 688
rect 1904 682 1912 683
rect 1924 688 1932 689
rect 1972 690 1980 691
rect 1924 683 1932 684
rect 1972 687 1980 688
rect 1924 680 1932 681
rect 1904 679 1912 680
rect 1972 682 1980 683
rect 1972 679 1980 680
rect 1924 666 1932 667
rect 1904 665 1912 666
rect 1904 662 1912 663
rect 1904 657 1912 658
rect 1924 663 1932 664
rect 1972 665 1980 666
rect 1924 658 1932 659
rect 1972 662 1980 663
rect 1924 655 1932 656
rect 1904 654 1912 655
rect 1972 657 1980 658
rect 1972 654 1980 655
rect 1924 641 1932 642
rect 1904 640 1912 641
rect 1904 637 1912 638
rect 1904 632 1912 633
rect 1924 638 1932 639
rect 1972 640 1980 641
rect 1924 633 1932 634
rect 1972 637 1980 638
rect 1924 630 1932 631
rect 1904 629 1912 630
rect 1972 632 1980 633
rect 1972 629 1980 630
rect 1924 616 1932 617
rect 1904 615 1912 616
rect 1904 612 1912 613
rect 1904 607 1912 608
rect 1924 613 1932 614
rect 1972 615 1980 616
rect 1924 608 1932 609
rect 1972 612 1980 613
rect 1924 605 1932 606
rect 1904 604 1912 605
rect 1972 607 1980 608
rect 1972 604 1980 605
rect 1924 591 1932 592
rect 1904 590 1912 591
rect 1904 587 1912 588
rect 1904 582 1912 583
rect 1924 588 1932 589
rect 1972 590 1980 591
rect 1924 583 1932 584
rect 1972 587 1980 588
rect 1924 580 1932 581
rect 1904 579 1912 580
rect 1972 582 1980 583
rect 1972 579 1980 580
rect 1924 566 1932 567
rect 1904 565 1912 566
rect 1904 562 1912 563
rect 1904 557 1912 558
rect 1924 563 1932 564
rect 1972 565 1980 566
rect 1924 558 1932 559
rect 1972 562 1980 563
rect 1924 555 1932 556
rect 1904 554 1912 555
rect 1972 557 1980 558
rect 1972 554 1980 555
rect 1924 541 1932 542
rect 1904 540 1912 541
rect 1904 537 1912 538
rect 1904 532 1912 533
rect 1924 538 1932 539
rect 1972 540 1980 541
rect 1924 533 1932 534
rect 1972 537 1980 538
rect 1924 530 1932 531
rect 1904 529 1912 530
rect 1972 532 1980 533
rect 1972 529 1980 530
rect 1924 516 1932 517
rect 1904 515 1912 516
rect 1904 512 1912 513
rect 1904 507 1912 508
rect 1924 513 1932 514
rect 1972 515 1980 516
rect 1924 508 1932 509
rect 1972 512 1980 513
rect 1924 505 1932 506
rect 1904 504 1912 505
rect 1972 507 1980 508
rect 1972 504 1980 505
rect 1924 491 1932 492
rect 1904 490 1912 491
rect 1904 487 1912 488
rect 1904 482 1912 483
rect 1924 488 1932 489
rect 1972 490 1980 491
rect 1924 483 1932 484
rect 1972 487 1980 488
rect 1924 480 1932 481
rect 1904 479 1912 480
rect 1972 482 1980 483
rect 1972 479 1980 480
rect 1924 466 1932 467
rect 1904 465 1912 466
rect 1904 462 1912 463
rect 1904 457 1912 458
rect 1924 463 1932 464
rect 1972 465 1980 466
rect 1924 458 1932 459
rect 1972 462 1980 463
rect 1924 455 1932 456
rect 1904 454 1912 455
rect 1972 457 1980 458
rect 1972 454 1980 455
rect 1924 441 1932 442
rect 1904 440 1912 441
rect 1904 437 1912 438
rect 1904 432 1912 433
rect 1924 438 1932 439
rect 1972 440 1980 441
rect 1924 433 1932 434
rect 1972 437 1980 438
rect 1924 430 1932 431
rect 1904 429 1912 430
rect 1972 432 1980 433
rect 1972 429 1980 430
rect 1924 416 1932 417
rect 1904 415 1912 416
rect 1904 412 1912 413
rect 1904 407 1912 408
rect 1924 413 1932 414
rect 1972 415 1980 416
rect 1924 408 1932 409
rect 1972 412 1980 413
rect 1924 405 1932 406
rect 1904 404 1912 405
rect 1972 407 1980 408
rect 1972 404 1980 405
rect 1924 391 1932 392
rect 1904 390 1912 391
rect 1904 387 1912 388
rect 1904 382 1912 383
rect 1924 388 1932 389
rect 1972 390 1980 391
rect 1924 383 1932 384
rect 1972 387 1980 388
rect 1924 380 1932 381
rect 1904 379 1912 380
rect 1972 382 1980 383
rect 1972 379 1980 380
rect 1924 366 1932 367
rect 1904 365 1912 366
rect 1904 362 1912 363
rect 1904 357 1912 358
rect 1924 363 1932 364
rect 1972 365 1980 366
rect 1924 358 1932 359
rect 1972 362 1980 363
rect 1924 355 1932 356
rect 1904 354 1912 355
rect 1972 357 1980 358
rect 1972 354 1980 355
rect 1924 341 1932 342
rect 1904 340 1912 341
rect 1904 337 1912 338
rect 1904 332 1912 333
rect 1924 338 1932 339
rect 1972 340 1980 341
rect 1924 333 1932 334
rect 1972 337 1980 338
rect 1924 330 1932 331
rect 1904 329 1912 330
rect 1972 332 1980 333
rect 1972 329 1980 330
rect 1924 316 1932 317
rect 1904 315 1912 316
rect 1904 312 1912 313
rect 1904 307 1912 308
rect 1924 313 1932 314
rect 1972 315 1980 316
rect 1924 308 1932 309
rect 1972 312 1980 313
rect 1924 305 1932 306
rect 1904 304 1912 305
rect 1972 307 1980 308
rect 1972 304 1980 305
rect 1924 291 1932 292
rect 1904 290 1912 291
rect 1904 287 1912 288
rect 1904 282 1912 283
rect 1924 288 1932 289
rect 1972 290 1980 291
rect 1924 283 1932 284
rect 1972 287 1980 288
rect 1924 280 1932 281
rect 1904 279 1912 280
rect 1972 282 1980 283
rect 1972 279 1980 280
rect 1924 266 1932 267
rect 1904 265 1912 266
rect 1904 262 1912 263
rect 1904 257 1912 258
rect 1924 263 1932 264
rect 1972 265 1980 266
rect 1924 258 1932 259
rect 1972 262 1980 263
rect 1924 255 1932 256
rect 1904 254 1912 255
rect 1972 257 1980 258
rect 1972 254 1980 255
rect 1924 241 1932 242
rect 1904 240 1912 241
rect 1904 237 1912 238
rect 1904 232 1912 233
rect 1924 238 1932 239
rect 1972 240 1980 241
rect 1924 233 1932 234
rect 1972 237 1980 238
rect 1924 230 1932 231
rect 1904 229 1912 230
rect 1972 232 1980 233
rect 1972 229 1980 230
rect 1924 216 1932 217
rect 1904 215 1912 216
rect 1904 212 1912 213
rect 1904 207 1912 208
rect 1924 213 1932 214
rect 1972 215 1980 216
rect 1924 208 1932 209
rect 1972 212 1980 213
rect 1924 205 1932 206
rect 1904 204 1912 205
rect 1972 207 1980 208
rect 1972 204 1980 205
rect 1924 191 1932 192
rect 1904 190 1912 191
rect 1904 187 1912 188
rect 1904 182 1912 183
rect 1924 188 1932 189
rect 1972 190 1980 191
rect 1924 183 1932 184
rect 1972 187 1980 188
rect 1924 180 1932 181
rect 1904 179 1912 180
rect 1972 182 1980 183
rect 1972 179 1980 180
rect 1924 166 1932 167
rect 1904 165 1912 166
rect 1904 162 1912 163
rect 1904 157 1912 158
rect 1924 163 1932 164
rect 1972 165 1980 166
rect 1924 158 1932 159
rect 1972 162 1980 163
rect 1924 155 1932 156
rect 1904 154 1912 155
rect 1972 157 1980 158
rect 1972 154 1980 155
rect 1924 141 1932 142
rect 1904 140 1912 141
rect 1904 137 1912 138
rect 1904 132 1912 133
rect 1924 138 1932 139
rect 1972 140 1980 141
rect 1924 133 1932 134
rect 1972 137 1980 138
rect 1924 130 1932 131
rect 1904 129 1912 130
rect 1972 132 1980 133
rect 1972 129 1980 130
rect 1924 116 1932 117
rect 1904 115 1912 116
rect 1904 112 1912 113
rect 1904 107 1912 108
rect 1924 113 1932 114
rect 1972 115 1980 116
rect 1924 108 1932 109
rect 1972 112 1980 113
rect 1924 105 1932 106
rect 1904 104 1912 105
rect 1972 107 1980 108
rect 1972 104 1980 105
rect 1924 91 1932 92
rect 1904 90 1912 91
rect 1904 87 1912 88
rect 1904 82 1912 83
rect 1924 88 1932 89
rect 1972 90 1980 91
rect 1924 83 1932 84
rect 1972 87 1980 88
rect 1924 80 1932 81
rect 1904 79 1912 80
rect 1972 82 1980 83
rect 1972 79 1980 80
rect 1924 66 1932 67
rect 1904 65 1912 66
rect 1904 62 1912 63
rect 1904 57 1912 58
rect 1924 63 1932 64
rect 1972 65 1980 66
rect 1924 58 1932 59
rect 1972 62 1980 63
rect 1924 55 1932 56
rect 1904 54 1912 55
rect 1972 57 1980 58
rect 1972 54 1980 55
rect 1924 41 1932 42
rect 1904 40 1912 41
rect 1904 37 1912 38
rect 1904 32 1912 33
rect 1924 38 1932 39
rect 1972 40 1980 41
rect 1924 33 1932 34
rect 1972 37 1980 38
rect 1924 30 1932 31
rect 1904 29 1912 30
rect 1972 32 1980 33
rect 1972 29 1980 30
<< metal1 >>
rect 1882 2026 1954 2029
rect 870 2018 1715 2026
rect 870 1888 878 2018
rect 928 2006 1704 2014
rect 20 1880 878 1888
rect 882 1984 998 2000
rect 1645 1984 1689 2000
rect 882 1876 916 1984
rect -36 1840 916 1876
rect 938 1910 1001 1926
rect -35 1778 5 1840
rect 43 1821 49 1828
rect 938 1823 976 1910
rect 1653 1889 1657 1897
rect 910 1807 976 1823
rect -34 1749 4 1778
rect -34 1733 30 1749
rect -34 1560 4 1733
rect 938 1725 976 1807
rect 1665 1799 1689 1984
rect 1642 1783 1689 1799
rect 1424 1742 1430 1751
rect 938 1709 1001 1725
rect 938 1675 976 1709
rect 909 1659 976 1675
rect 915 1635 920 1643
rect 910 1617 917 1623
rect 938 1577 976 1659
rect 1424 1663 1430 1664
rect 1665 1651 1689 1783
rect 1642 1635 1689 1651
rect 938 1561 1000 1577
rect 1096 1561 1229 1566
rect -34 1544 30 1560
rect 938 1554 1653 1561
rect -34 1359 4 1544
rect 938 1538 1002 1554
rect 1096 1545 1229 1554
rect 910 1446 929 1454
rect 938 1433 976 1538
rect 1336 1477 1344 1494
rect 1665 1480 1689 1635
rect 1642 1464 1647 1480
rect 1654 1464 1689 1480
rect 910 1417 976 1433
rect 938 1406 976 1417
rect 1675 1418 1689 1464
rect 1696 1431 1704 2006
rect 1707 1442 1715 2018
rect 1796 2019 1867 2026
rect 1796 1431 1804 2019
rect 1696 1423 1804 1431
rect 1675 1414 1711 1418
rect 1750 1414 1770 1418
rect 938 1390 999 1406
rect 1655 1390 1670 1406
rect 1682 1398 1707 1411
rect -34 1339 30 1359
rect -34 1124 4 1339
rect 938 1229 976 1390
rect 1661 1381 1688 1390
rect 1699 1387 1707 1398
rect 1752 1410 1756 1414
rect 1699 1383 1711 1387
rect 1424 1372 1433 1375
rect 1427 1371 1433 1372
rect 1671 1363 1680 1372
rect 1684 1366 1688 1381
rect 1762 1380 1766 1390
rect 1796 1387 1804 1423
rect 1792 1383 1804 1387
rect 1766 1370 1785 1373
rect 1752 1366 1756 1370
rect 1763 1369 1785 1370
rect 1684 1362 1712 1366
rect 1750 1362 1770 1366
rect 1796 1363 1804 1383
rect 1778 1358 1804 1363
rect 1778 1348 1785 1358
rect 1796 1348 1804 1358
rect 1882 2014 1886 2026
rect 1894 2016 1904 2020
rect 1886 2008 1890 2012
rect 1897 2010 1901 2016
rect 1916 2015 1920 2023
rect 1932 2019 1935 2021
rect 1939 2019 1942 2021
rect 1932 2018 1942 2019
rect 1950 2015 1954 2026
rect 1962 2016 1972 2020
rect 1912 2008 1916 2012
rect 1920 2009 1924 2013
rect 1882 1989 1886 2006
rect 1894 2002 1904 2003
rect 1894 2000 1897 2002
rect 1901 2000 1904 2002
rect 1894 1991 1904 1995
rect 1886 1983 1890 1987
rect 1897 1985 1901 1991
rect 1916 1990 1920 2006
rect 1935 2005 1939 2011
rect 1946 2009 1950 2013
rect 1954 2008 1958 2012
rect 1965 2010 1969 2016
rect 1984 2015 1988 2023
rect 1980 2008 1984 2012
rect 1932 2001 1942 2005
rect 1932 1994 1935 1996
rect 1939 1994 1942 1996
rect 1932 1993 1942 1994
rect 1950 1990 1954 2006
rect 1962 2002 1972 2003
rect 1962 2000 1965 2002
rect 1969 2000 1972 2002
rect 1962 1991 1972 1995
rect 1912 1983 1916 1987
rect 1920 1984 1924 1988
rect 1882 1964 1886 1981
rect 1894 1977 1904 1978
rect 1894 1975 1897 1977
rect 1901 1975 1904 1977
rect 1894 1966 1904 1970
rect 1886 1958 1890 1962
rect 1897 1960 1901 1966
rect 1916 1965 1920 1981
rect 1935 1980 1939 1986
rect 1946 1984 1950 1988
rect 1954 1983 1958 1987
rect 1965 1985 1969 1991
rect 1984 1990 1988 2006
rect 1980 1983 1984 1987
rect 1932 1976 1942 1980
rect 1932 1969 1935 1971
rect 1939 1969 1942 1971
rect 1932 1968 1942 1969
rect 1950 1965 1954 1981
rect 1962 1977 1972 1978
rect 1962 1975 1965 1977
rect 1969 1975 1972 1977
rect 1962 1966 1972 1970
rect 1912 1958 1916 1962
rect 1920 1959 1924 1963
rect 1882 1939 1886 1956
rect 1894 1952 1904 1953
rect 1894 1950 1897 1952
rect 1901 1950 1904 1952
rect 1894 1941 1904 1945
rect 1886 1933 1890 1937
rect 1897 1935 1901 1941
rect 1916 1940 1920 1956
rect 1935 1955 1939 1961
rect 1946 1959 1950 1963
rect 1954 1958 1958 1962
rect 1965 1960 1969 1966
rect 1984 1965 1988 1981
rect 1980 1958 1984 1962
rect 1932 1951 1942 1955
rect 1932 1944 1935 1946
rect 1939 1944 1942 1946
rect 1932 1943 1942 1944
rect 1950 1940 1954 1956
rect 1962 1952 1972 1953
rect 1962 1950 1965 1952
rect 1969 1950 1972 1952
rect 1962 1941 1972 1945
rect 1912 1933 1916 1937
rect 1920 1934 1924 1938
rect 1882 1914 1886 1931
rect 1894 1927 1904 1928
rect 1894 1925 1897 1927
rect 1901 1925 1904 1927
rect 1894 1916 1904 1920
rect 1886 1908 1890 1912
rect 1897 1910 1901 1916
rect 1916 1915 1920 1931
rect 1935 1930 1939 1936
rect 1946 1934 1950 1938
rect 1954 1933 1958 1937
rect 1965 1935 1969 1941
rect 1984 1940 1988 1956
rect 1980 1933 1984 1937
rect 1932 1926 1942 1930
rect 1932 1919 1935 1921
rect 1939 1919 1942 1921
rect 1932 1918 1942 1919
rect 1950 1915 1954 1931
rect 1962 1927 1972 1928
rect 1962 1925 1965 1927
rect 1969 1925 1972 1927
rect 1962 1916 1972 1920
rect 1912 1908 1916 1912
rect 1920 1909 1924 1913
rect 1882 1889 1886 1906
rect 1894 1902 1904 1903
rect 1894 1900 1897 1902
rect 1901 1900 1904 1902
rect 1894 1891 1904 1895
rect 1886 1883 1890 1887
rect 1897 1885 1901 1891
rect 1916 1890 1920 1906
rect 1935 1905 1939 1911
rect 1946 1909 1950 1913
rect 1954 1908 1958 1912
rect 1965 1910 1969 1916
rect 1984 1915 1988 1931
rect 1980 1908 1984 1912
rect 1932 1901 1942 1905
rect 1932 1894 1935 1896
rect 1939 1894 1942 1896
rect 1932 1893 1942 1894
rect 1950 1890 1954 1906
rect 1962 1902 1972 1903
rect 1962 1900 1965 1902
rect 1969 1900 1972 1902
rect 1962 1891 1972 1895
rect 1912 1883 1916 1887
rect 1920 1884 1924 1888
rect 1882 1864 1886 1881
rect 1894 1877 1904 1878
rect 1894 1875 1897 1877
rect 1901 1875 1904 1877
rect 1894 1866 1904 1870
rect 1886 1858 1890 1862
rect 1897 1860 1901 1866
rect 1916 1865 1920 1881
rect 1935 1880 1939 1886
rect 1946 1884 1950 1888
rect 1954 1883 1958 1887
rect 1965 1885 1969 1891
rect 1984 1890 1988 1906
rect 1980 1883 1984 1887
rect 1932 1876 1942 1880
rect 1932 1869 1935 1871
rect 1939 1869 1942 1871
rect 1932 1868 1942 1869
rect 1950 1865 1954 1881
rect 1962 1877 1972 1878
rect 1962 1875 1965 1877
rect 1969 1875 1972 1877
rect 1962 1866 1972 1870
rect 1912 1858 1916 1862
rect 1920 1859 1924 1863
rect 1882 1839 1886 1856
rect 1894 1852 1904 1853
rect 1894 1850 1897 1852
rect 1901 1850 1904 1852
rect 1894 1841 1904 1845
rect 1886 1833 1890 1837
rect 1897 1835 1901 1841
rect 1916 1840 1920 1856
rect 1935 1855 1939 1861
rect 1946 1859 1950 1863
rect 1954 1858 1958 1862
rect 1965 1860 1969 1866
rect 1984 1865 1988 1881
rect 1980 1858 1984 1862
rect 1932 1851 1942 1855
rect 1932 1844 1935 1846
rect 1939 1844 1942 1846
rect 1932 1843 1942 1844
rect 1950 1840 1954 1856
rect 1962 1852 1972 1853
rect 1962 1850 1965 1852
rect 1969 1850 1972 1852
rect 1962 1841 1972 1845
rect 1912 1833 1916 1837
rect 1920 1834 1924 1838
rect 1882 1814 1886 1831
rect 1894 1827 1904 1828
rect 1894 1825 1897 1827
rect 1901 1825 1904 1827
rect 1894 1816 1904 1820
rect 1886 1808 1890 1812
rect 1897 1810 1901 1816
rect 1916 1815 1920 1831
rect 1935 1830 1939 1836
rect 1946 1834 1950 1838
rect 1954 1833 1958 1837
rect 1965 1835 1969 1841
rect 1984 1840 1988 1856
rect 1980 1833 1984 1837
rect 1932 1826 1942 1830
rect 1932 1819 1935 1821
rect 1939 1819 1942 1821
rect 1932 1818 1942 1819
rect 1950 1815 1954 1831
rect 1962 1827 1972 1828
rect 1962 1825 1965 1827
rect 1969 1825 1972 1827
rect 1962 1816 1972 1820
rect 1912 1808 1916 1812
rect 1920 1809 1924 1813
rect 1882 1789 1886 1806
rect 1894 1802 1904 1803
rect 1894 1800 1897 1802
rect 1901 1800 1904 1802
rect 1894 1791 1904 1795
rect 1886 1783 1890 1787
rect 1897 1785 1901 1791
rect 1916 1790 1920 1806
rect 1935 1805 1939 1811
rect 1946 1809 1950 1813
rect 1954 1808 1958 1812
rect 1965 1810 1969 1816
rect 1984 1815 1988 1831
rect 1980 1808 1984 1812
rect 1932 1801 1942 1805
rect 1932 1794 1935 1796
rect 1939 1794 1942 1796
rect 1932 1793 1942 1794
rect 1950 1790 1954 1806
rect 1962 1802 1972 1803
rect 1962 1800 1965 1802
rect 1969 1800 1972 1802
rect 1962 1791 1972 1795
rect 1912 1783 1916 1787
rect 1920 1784 1924 1788
rect 1882 1764 1886 1781
rect 1894 1777 1904 1778
rect 1894 1775 1897 1777
rect 1901 1775 1904 1777
rect 1894 1766 1904 1770
rect 1886 1758 1890 1762
rect 1897 1760 1901 1766
rect 1916 1765 1920 1781
rect 1935 1780 1939 1786
rect 1946 1784 1950 1788
rect 1954 1783 1958 1787
rect 1965 1785 1969 1791
rect 1984 1790 1988 1806
rect 1980 1783 1984 1787
rect 1932 1776 1942 1780
rect 1932 1769 1935 1771
rect 1939 1769 1942 1771
rect 1932 1768 1942 1769
rect 1950 1765 1954 1781
rect 1962 1777 1972 1778
rect 1962 1775 1965 1777
rect 1969 1775 1972 1777
rect 1962 1766 1972 1770
rect 1912 1758 1916 1762
rect 1920 1759 1924 1763
rect 1882 1739 1886 1756
rect 1894 1752 1904 1753
rect 1894 1750 1897 1752
rect 1901 1750 1904 1752
rect 1894 1741 1904 1745
rect 1886 1733 1890 1737
rect 1897 1735 1901 1741
rect 1916 1740 1920 1756
rect 1935 1755 1939 1761
rect 1946 1759 1950 1763
rect 1954 1758 1958 1762
rect 1965 1760 1969 1766
rect 1984 1765 1988 1781
rect 1980 1758 1984 1762
rect 1932 1751 1942 1755
rect 1932 1744 1935 1746
rect 1939 1744 1942 1746
rect 1932 1743 1942 1744
rect 1950 1740 1954 1756
rect 1962 1752 1972 1753
rect 1962 1750 1965 1752
rect 1969 1750 1972 1752
rect 1962 1741 1972 1745
rect 1912 1733 1916 1737
rect 1920 1734 1924 1738
rect 1882 1714 1886 1731
rect 1894 1727 1904 1728
rect 1894 1725 1897 1727
rect 1901 1725 1904 1727
rect 1894 1716 1904 1720
rect 1886 1708 1890 1712
rect 1897 1710 1901 1716
rect 1916 1715 1920 1731
rect 1935 1730 1939 1736
rect 1946 1734 1950 1738
rect 1954 1733 1958 1737
rect 1965 1735 1969 1741
rect 1984 1740 1988 1756
rect 1980 1733 1984 1737
rect 1932 1726 1942 1730
rect 1932 1719 1935 1721
rect 1939 1719 1942 1721
rect 1932 1718 1942 1719
rect 1950 1715 1954 1731
rect 1962 1727 1972 1728
rect 1962 1725 1965 1727
rect 1969 1725 1972 1727
rect 1962 1716 1972 1720
rect 1912 1708 1916 1712
rect 1920 1709 1924 1713
rect 1882 1689 1886 1706
rect 1894 1702 1904 1703
rect 1894 1700 1897 1702
rect 1901 1700 1904 1702
rect 1894 1691 1904 1695
rect 1886 1683 1890 1687
rect 1897 1685 1901 1691
rect 1916 1690 1920 1706
rect 1935 1705 1939 1711
rect 1946 1709 1950 1713
rect 1954 1708 1958 1712
rect 1965 1710 1969 1716
rect 1984 1715 1988 1731
rect 1980 1708 1984 1712
rect 1932 1701 1942 1705
rect 1932 1694 1935 1696
rect 1939 1694 1942 1696
rect 1932 1693 1942 1694
rect 1950 1690 1954 1706
rect 1962 1702 1972 1703
rect 1962 1700 1965 1702
rect 1969 1700 1972 1702
rect 1962 1691 1972 1695
rect 1912 1683 1916 1687
rect 1920 1684 1924 1688
rect 1882 1664 1886 1681
rect 1894 1677 1904 1678
rect 1894 1675 1897 1677
rect 1901 1675 1904 1677
rect 1894 1666 1904 1670
rect 1886 1658 1890 1662
rect 1897 1660 1901 1666
rect 1916 1665 1920 1681
rect 1935 1680 1939 1686
rect 1946 1684 1950 1688
rect 1954 1683 1958 1687
rect 1965 1685 1969 1691
rect 1984 1690 1988 1706
rect 1980 1683 1984 1687
rect 1932 1676 1942 1680
rect 1932 1669 1935 1671
rect 1939 1669 1942 1671
rect 1932 1668 1942 1669
rect 1950 1665 1954 1681
rect 1962 1677 1972 1678
rect 1962 1675 1965 1677
rect 1969 1675 1972 1677
rect 1962 1666 1972 1670
rect 1912 1658 1916 1662
rect 1920 1659 1924 1663
rect 1882 1639 1886 1656
rect 1894 1652 1904 1653
rect 1894 1650 1897 1652
rect 1901 1650 1904 1652
rect 1894 1641 1904 1645
rect 1886 1633 1890 1637
rect 1897 1635 1901 1641
rect 1916 1640 1920 1656
rect 1935 1655 1939 1661
rect 1946 1659 1950 1663
rect 1954 1658 1958 1662
rect 1965 1660 1969 1666
rect 1984 1665 1988 1681
rect 1980 1658 1984 1662
rect 1932 1651 1942 1655
rect 1932 1644 1935 1646
rect 1939 1644 1942 1646
rect 1932 1643 1942 1644
rect 1950 1640 1954 1656
rect 1962 1652 1972 1653
rect 1962 1650 1965 1652
rect 1969 1650 1972 1652
rect 1962 1641 1972 1645
rect 1912 1633 1916 1637
rect 1920 1634 1924 1638
rect 1882 1614 1886 1631
rect 1894 1627 1904 1628
rect 1894 1625 1897 1627
rect 1901 1625 1904 1627
rect 1894 1616 1904 1620
rect 1886 1608 1890 1612
rect 1897 1610 1901 1616
rect 1916 1615 1920 1631
rect 1935 1630 1939 1636
rect 1946 1634 1950 1638
rect 1954 1633 1958 1637
rect 1965 1635 1969 1641
rect 1984 1640 1988 1656
rect 1980 1633 1984 1637
rect 1932 1626 1942 1630
rect 1932 1619 1935 1621
rect 1939 1619 1942 1621
rect 1932 1618 1942 1619
rect 1950 1615 1954 1631
rect 1962 1627 1972 1628
rect 1962 1625 1965 1627
rect 1969 1625 1972 1627
rect 1962 1616 1972 1620
rect 1912 1608 1916 1612
rect 1920 1609 1924 1613
rect 1882 1589 1886 1606
rect 1894 1602 1904 1603
rect 1894 1600 1897 1602
rect 1901 1600 1904 1602
rect 1894 1591 1904 1595
rect 1886 1583 1890 1587
rect 1897 1585 1901 1591
rect 1916 1590 1920 1606
rect 1935 1605 1939 1611
rect 1946 1609 1950 1613
rect 1954 1608 1958 1612
rect 1965 1610 1969 1616
rect 1984 1615 1988 1631
rect 1980 1608 1984 1612
rect 1932 1601 1942 1605
rect 1932 1594 1935 1596
rect 1939 1594 1942 1596
rect 1932 1593 1942 1594
rect 1950 1590 1954 1606
rect 1962 1602 1972 1603
rect 1962 1600 1965 1602
rect 1969 1600 1972 1602
rect 1962 1591 1972 1595
rect 1912 1583 1916 1587
rect 1920 1584 1924 1588
rect 1882 1564 1886 1581
rect 1894 1577 1904 1578
rect 1894 1575 1897 1577
rect 1901 1575 1904 1577
rect 1894 1566 1904 1570
rect 1886 1558 1890 1562
rect 1897 1560 1901 1566
rect 1916 1565 1920 1581
rect 1935 1580 1939 1586
rect 1946 1584 1950 1588
rect 1954 1583 1958 1587
rect 1965 1585 1969 1591
rect 1984 1590 1988 1606
rect 1980 1583 1984 1587
rect 1932 1576 1942 1580
rect 1932 1569 1935 1571
rect 1939 1569 1942 1571
rect 1932 1568 1942 1569
rect 1950 1565 1954 1581
rect 1962 1577 1972 1578
rect 1962 1575 1965 1577
rect 1969 1575 1972 1577
rect 1962 1566 1972 1570
rect 1912 1558 1916 1562
rect 1920 1559 1924 1563
rect 1882 1539 1886 1556
rect 1894 1552 1904 1553
rect 1894 1550 1897 1552
rect 1901 1550 1904 1552
rect 1894 1541 1904 1545
rect 1886 1533 1890 1537
rect 1897 1535 1901 1541
rect 1916 1540 1920 1556
rect 1935 1555 1939 1561
rect 1946 1559 1950 1563
rect 1954 1558 1958 1562
rect 1965 1560 1969 1566
rect 1984 1565 1988 1581
rect 1980 1558 1984 1562
rect 1932 1551 1942 1555
rect 1932 1544 1935 1546
rect 1939 1544 1942 1546
rect 1932 1543 1942 1544
rect 1950 1540 1954 1556
rect 1962 1552 1972 1553
rect 1962 1550 1965 1552
rect 1969 1550 1972 1552
rect 1962 1541 1972 1545
rect 1912 1533 1916 1537
rect 1920 1534 1924 1538
rect 1882 1514 1886 1531
rect 1894 1527 1904 1528
rect 1894 1525 1897 1527
rect 1901 1525 1904 1527
rect 1894 1516 1904 1520
rect 1886 1508 1890 1512
rect 1897 1510 1901 1516
rect 1916 1515 1920 1531
rect 1935 1530 1939 1536
rect 1946 1534 1950 1538
rect 1954 1533 1958 1537
rect 1965 1535 1969 1541
rect 1984 1540 1988 1556
rect 1980 1533 1984 1537
rect 1932 1526 1942 1530
rect 1932 1519 1935 1521
rect 1939 1519 1942 1521
rect 1932 1518 1942 1519
rect 1950 1515 1954 1531
rect 1962 1527 1972 1528
rect 1962 1525 1965 1527
rect 1969 1525 1972 1527
rect 1962 1516 1972 1520
rect 1912 1508 1916 1512
rect 1920 1509 1924 1513
rect 1882 1489 1886 1506
rect 1894 1502 1904 1503
rect 1894 1500 1897 1502
rect 1901 1500 1904 1502
rect 1894 1491 1904 1495
rect 1886 1483 1890 1487
rect 1897 1485 1901 1491
rect 1916 1490 1920 1506
rect 1935 1505 1939 1511
rect 1946 1509 1950 1513
rect 1954 1508 1958 1512
rect 1965 1510 1969 1516
rect 1984 1515 1988 1531
rect 1980 1508 1984 1512
rect 1932 1501 1942 1505
rect 1932 1494 1935 1496
rect 1939 1494 1942 1496
rect 1932 1493 1942 1494
rect 1950 1490 1954 1506
rect 1962 1502 1972 1503
rect 1962 1500 1965 1502
rect 1969 1500 1972 1502
rect 1962 1491 1972 1495
rect 1912 1483 1916 1487
rect 1920 1484 1924 1488
rect 1882 1464 1886 1481
rect 1894 1477 1904 1478
rect 1894 1475 1897 1477
rect 1901 1475 1904 1477
rect 1894 1466 1904 1470
rect 1886 1458 1890 1462
rect 1897 1460 1901 1466
rect 1916 1465 1920 1481
rect 1935 1480 1939 1486
rect 1946 1484 1950 1488
rect 1954 1483 1958 1487
rect 1965 1485 1969 1491
rect 1984 1490 1988 1506
rect 1980 1483 1984 1487
rect 1932 1476 1942 1480
rect 1932 1469 1935 1471
rect 1939 1469 1942 1471
rect 1932 1468 1942 1469
rect 1950 1465 1954 1481
rect 1962 1477 1972 1478
rect 1962 1475 1965 1477
rect 1969 1475 1972 1477
rect 1962 1466 1972 1470
rect 1912 1458 1916 1462
rect 1920 1459 1924 1463
rect 1882 1439 1886 1456
rect 1894 1452 1904 1453
rect 1894 1450 1897 1452
rect 1901 1450 1904 1452
rect 1894 1441 1904 1445
rect 1886 1433 1890 1437
rect 1897 1435 1901 1441
rect 1916 1440 1920 1456
rect 1935 1455 1939 1461
rect 1946 1459 1950 1463
rect 1954 1458 1958 1462
rect 1965 1460 1969 1466
rect 1984 1465 1988 1481
rect 1980 1458 1984 1462
rect 1932 1451 1942 1455
rect 1932 1444 1935 1446
rect 1939 1444 1942 1446
rect 1932 1443 1942 1444
rect 1950 1440 1954 1456
rect 1962 1452 1972 1453
rect 1962 1450 1965 1452
rect 1969 1450 1972 1452
rect 1962 1441 1972 1445
rect 1912 1433 1916 1437
rect 1920 1434 1924 1438
rect 1882 1414 1886 1431
rect 1894 1427 1904 1428
rect 1894 1425 1897 1427
rect 1901 1425 1904 1427
rect 1894 1416 1904 1420
rect 1886 1408 1890 1412
rect 1897 1410 1901 1416
rect 1916 1415 1920 1431
rect 1935 1430 1939 1436
rect 1946 1434 1950 1438
rect 1954 1433 1958 1437
rect 1965 1435 1969 1441
rect 1984 1440 1988 1456
rect 1980 1433 1984 1437
rect 1932 1426 1942 1430
rect 1932 1419 1935 1421
rect 1939 1419 1942 1421
rect 1932 1418 1942 1419
rect 1950 1415 1954 1431
rect 1962 1427 1972 1428
rect 1962 1425 1965 1427
rect 1969 1425 1972 1427
rect 1962 1416 1972 1420
rect 1912 1408 1916 1412
rect 1920 1409 1924 1413
rect 1882 1389 1886 1406
rect 1894 1402 1904 1403
rect 1894 1400 1897 1402
rect 1901 1400 1904 1402
rect 1894 1391 1904 1395
rect 1886 1383 1890 1387
rect 1897 1385 1901 1391
rect 1916 1390 1920 1406
rect 1935 1405 1939 1411
rect 1946 1409 1950 1413
rect 1954 1408 1958 1412
rect 1965 1410 1969 1416
rect 1984 1415 1988 1431
rect 1980 1408 1984 1412
rect 1932 1401 1942 1405
rect 1932 1394 1935 1396
rect 1939 1394 1942 1396
rect 1932 1393 1942 1394
rect 1950 1390 1954 1406
rect 1962 1402 1972 1403
rect 1962 1400 1965 1402
rect 1969 1400 1972 1402
rect 1962 1391 1972 1395
rect 1912 1383 1916 1387
rect 1920 1384 1924 1388
rect 1882 1364 1886 1381
rect 1894 1377 1904 1378
rect 1894 1375 1897 1377
rect 1901 1375 1904 1377
rect 1894 1366 1904 1370
rect 1886 1358 1890 1362
rect 1897 1360 1901 1366
rect 1916 1365 1920 1381
rect 1935 1380 1939 1386
rect 1946 1384 1950 1388
rect 1954 1383 1958 1387
rect 1965 1385 1969 1391
rect 1984 1390 1988 1406
rect 1980 1383 1984 1387
rect 1932 1376 1942 1380
rect 1932 1369 1935 1371
rect 1939 1369 1942 1371
rect 1932 1368 1942 1369
rect 1950 1365 1954 1381
rect 1962 1377 1972 1378
rect 1962 1375 1965 1377
rect 1969 1375 1972 1377
rect 1962 1366 1972 1370
rect 1912 1358 1916 1362
rect 1920 1359 1924 1363
rect 1775 1314 1824 1318
rect 1775 1291 1793 1295
rect 1779 1260 1786 1264
rect 910 1221 976 1229
rect 916 1198 920 1221
rect 938 1205 976 1221
rect 991 1218 999 1226
rect 938 1189 998 1205
rect 1778 1189 1782 1193
rect 906 1178 910 1188
rect 918 1181 921 1185
rect 916 1124 920 1158
rect -34 1116 30 1124
rect 907 1116 920 1124
rect -34 893 4 1116
rect 20 1022 48 1039
rect 938 1021 976 1189
rect 1743 1115 1746 1116
rect 1743 1100 1747 1115
rect 1739 1096 1747 1100
rect 1750 1101 1754 1105
rect 1739 1093 1743 1096
rect 1757 1093 1761 1117
rect 1768 1097 1772 1101
rect 1729 1065 1733 1075
rect 1747 1072 1751 1075
rect 1767 1072 1771 1075
rect 1740 1068 1771 1072
rect 1747 1065 1751 1068
rect 987 1049 1513 1052
rect 1729 1049 1733 1055
rect 987 1044 1733 1049
rect 1739 1044 1743 1055
rect 1767 1044 1771 1055
rect 1739 1040 1771 1044
rect 987 1028 1744 1036
rect 1755 1021 1759 1040
rect 1782 1036 1786 1189
rect 1789 1101 1793 1291
rect 1770 1028 1786 1036
rect 1796 1028 1800 1256
rect 1804 1028 1808 1264
rect 1812 1028 1816 1158
rect 1820 1028 1824 1314
rect 1828 1028 1836 1105
rect 1844 1028 1852 1344
rect 1882 1339 1886 1356
rect 1894 1352 1904 1353
rect 1894 1350 1897 1352
rect 1901 1350 1904 1352
rect 1894 1341 1904 1345
rect 1886 1333 1890 1337
rect 1897 1335 1901 1341
rect 1916 1340 1920 1356
rect 1935 1355 1939 1361
rect 1946 1359 1950 1363
rect 1954 1358 1958 1362
rect 1965 1360 1969 1366
rect 1984 1365 1988 1381
rect 1980 1358 1984 1362
rect 1932 1351 1942 1355
rect 1932 1344 1935 1346
rect 1939 1344 1942 1346
rect 1932 1343 1942 1344
rect 1950 1340 1954 1356
rect 1962 1352 1972 1353
rect 1962 1350 1965 1352
rect 1969 1350 1972 1352
rect 1962 1341 1972 1345
rect 1912 1333 1916 1337
rect 1920 1334 1924 1338
rect 1882 1314 1886 1331
rect 1894 1327 1904 1328
rect 1894 1325 1897 1327
rect 1901 1325 1904 1327
rect 1894 1316 1904 1320
rect 1886 1308 1890 1312
rect 1897 1310 1901 1316
rect 1916 1315 1920 1331
rect 1935 1330 1939 1336
rect 1946 1334 1950 1338
rect 1954 1333 1958 1337
rect 1965 1335 1969 1341
rect 1984 1340 1988 1356
rect 1980 1333 1984 1337
rect 1932 1326 1942 1330
rect 1932 1319 1935 1321
rect 1939 1319 1942 1321
rect 1932 1318 1942 1319
rect 1950 1315 1954 1331
rect 1962 1327 1972 1328
rect 1962 1325 1965 1327
rect 1969 1325 1972 1327
rect 1962 1316 1972 1320
rect 1912 1308 1916 1312
rect 1920 1309 1924 1313
rect 1882 1289 1886 1306
rect 1894 1302 1904 1303
rect 1894 1300 1897 1302
rect 1901 1300 1904 1302
rect 1894 1291 1904 1295
rect 1886 1283 1890 1287
rect 1897 1285 1901 1291
rect 1916 1290 1920 1306
rect 1935 1305 1939 1311
rect 1946 1309 1950 1313
rect 1954 1308 1958 1312
rect 1965 1310 1969 1316
rect 1984 1315 1988 1331
rect 1980 1308 1984 1312
rect 1932 1301 1942 1305
rect 1932 1294 1935 1296
rect 1939 1294 1942 1296
rect 1932 1293 1942 1294
rect 1950 1290 1954 1306
rect 1962 1302 1972 1303
rect 1962 1300 1965 1302
rect 1969 1300 1972 1302
rect 1962 1291 1972 1295
rect 1912 1283 1916 1287
rect 1920 1284 1924 1288
rect 1882 1264 1886 1281
rect 1894 1277 1904 1278
rect 1894 1275 1897 1277
rect 1901 1275 1904 1277
rect 1894 1266 1904 1270
rect 1886 1258 1890 1262
rect 1897 1260 1901 1266
rect 1916 1265 1920 1281
rect 1935 1280 1939 1286
rect 1946 1284 1950 1288
rect 1954 1283 1958 1287
rect 1965 1285 1969 1291
rect 1984 1290 1988 1306
rect 1980 1283 1984 1287
rect 1932 1276 1942 1280
rect 1932 1269 1935 1271
rect 1939 1269 1942 1271
rect 1932 1268 1942 1269
rect 1950 1265 1954 1281
rect 1962 1277 1972 1278
rect 1962 1275 1965 1277
rect 1969 1275 1972 1277
rect 1962 1266 1972 1270
rect 1912 1258 1916 1262
rect 1920 1259 1924 1263
rect 1882 1239 1886 1256
rect 1894 1252 1904 1253
rect 1894 1250 1897 1252
rect 1901 1250 1904 1252
rect 1894 1241 1904 1245
rect 1886 1233 1890 1237
rect 1897 1235 1901 1241
rect 1916 1240 1920 1256
rect 1935 1255 1939 1261
rect 1946 1259 1950 1263
rect 1954 1258 1958 1262
rect 1965 1260 1969 1266
rect 1984 1265 1988 1281
rect 1980 1258 1984 1262
rect 1932 1251 1942 1255
rect 1932 1244 1935 1246
rect 1939 1244 1942 1246
rect 1932 1243 1942 1244
rect 1950 1240 1954 1256
rect 1962 1252 1972 1253
rect 1962 1250 1965 1252
rect 1969 1250 1972 1252
rect 1962 1241 1972 1245
rect 1912 1233 1916 1237
rect 1920 1234 1924 1238
rect 1882 1214 1886 1231
rect 1894 1227 1904 1228
rect 1894 1225 1897 1227
rect 1901 1225 1904 1227
rect 1894 1216 1904 1220
rect 1886 1208 1890 1212
rect 1897 1210 1901 1216
rect 1916 1215 1920 1231
rect 1935 1230 1939 1236
rect 1946 1234 1950 1238
rect 1954 1233 1958 1237
rect 1965 1235 1969 1241
rect 1984 1240 1988 1256
rect 1980 1233 1984 1237
rect 1932 1226 1942 1230
rect 1932 1219 1935 1221
rect 1939 1219 1942 1221
rect 1932 1218 1942 1219
rect 1950 1215 1954 1231
rect 1962 1227 1972 1228
rect 1962 1225 1965 1227
rect 1969 1225 1972 1227
rect 1962 1216 1972 1220
rect 1912 1208 1916 1212
rect 1920 1209 1924 1213
rect 1882 1189 1886 1206
rect 1894 1202 1904 1203
rect 1894 1200 1897 1202
rect 1901 1200 1904 1202
rect 1894 1191 1904 1195
rect 1886 1183 1890 1187
rect 1897 1185 1901 1191
rect 1916 1190 1920 1206
rect 1935 1205 1939 1211
rect 1946 1209 1950 1213
rect 1954 1208 1958 1212
rect 1965 1210 1969 1216
rect 1984 1215 1988 1231
rect 1980 1208 1984 1212
rect 1932 1201 1942 1205
rect 1932 1194 1935 1196
rect 1939 1194 1942 1196
rect 1932 1193 1942 1194
rect 1950 1190 1954 1206
rect 1962 1202 1972 1203
rect 1962 1200 1965 1202
rect 1969 1200 1972 1202
rect 1962 1191 1972 1195
rect 1912 1183 1916 1187
rect 1920 1184 1924 1188
rect 1882 1164 1886 1181
rect 1894 1177 1904 1178
rect 1894 1175 1897 1177
rect 1901 1175 1904 1177
rect 1894 1166 1904 1170
rect 1886 1158 1890 1162
rect 1897 1160 1901 1166
rect 1916 1165 1920 1181
rect 1935 1180 1939 1186
rect 1946 1184 1950 1188
rect 1954 1183 1958 1187
rect 1965 1185 1969 1191
rect 1984 1190 1988 1206
rect 1980 1183 1984 1187
rect 1932 1176 1942 1180
rect 1932 1169 1935 1171
rect 1939 1169 1942 1171
rect 1932 1168 1942 1169
rect 1950 1165 1954 1181
rect 1962 1177 1972 1178
rect 1962 1175 1965 1177
rect 1969 1175 1972 1177
rect 1962 1166 1972 1170
rect 1912 1158 1916 1162
rect 1920 1159 1924 1163
rect 1882 1139 1886 1156
rect 1894 1152 1904 1153
rect 1894 1150 1897 1152
rect 1901 1150 1904 1152
rect 1894 1141 1904 1145
rect 1886 1133 1890 1137
rect 1897 1135 1901 1141
rect 1916 1140 1920 1156
rect 1935 1155 1939 1161
rect 1946 1159 1950 1163
rect 1954 1158 1958 1162
rect 1965 1160 1969 1166
rect 1984 1165 1988 1181
rect 1980 1158 1984 1162
rect 1932 1151 1942 1155
rect 1932 1144 1935 1146
rect 1939 1144 1942 1146
rect 1932 1143 1942 1144
rect 1950 1140 1954 1156
rect 1962 1152 1972 1153
rect 1962 1150 1965 1152
rect 1969 1150 1972 1152
rect 1962 1141 1972 1145
rect 1912 1133 1916 1137
rect 1920 1134 1924 1138
rect 1882 1114 1886 1131
rect 1894 1127 1904 1128
rect 1894 1125 1897 1127
rect 1901 1125 1904 1127
rect 1894 1116 1904 1120
rect 1886 1108 1890 1112
rect 1897 1110 1901 1116
rect 1916 1115 1920 1131
rect 1935 1130 1939 1136
rect 1946 1134 1950 1138
rect 1954 1133 1958 1137
rect 1965 1135 1969 1141
rect 1984 1140 1988 1156
rect 1980 1133 1984 1137
rect 1932 1126 1942 1130
rect 1932 1119 1935 1121
rect 1939 1119 1942 1121
rect 1932 1118 1942 1119
rect 1950 1115 1954 1131
rect 1962 1127 1972 1128
rect 1962 1125 1965 1127
rect 1969 1125 1972 1127
rect 1962 1116 1972 1120
rect 1912 1108 1916 1112
rect 1920 1109 1924 1113
rect 1882 1089 1886 1106
rect 1894 1102 1904 1103
rect 1894 1100 1897 1102
rect 1901 1100 1904 1102
rect 1894 1091 1904 1095
rect 1886 1083 1890 1087
rect 1897 1085 1901 1091
rect 1916 1090 1920 1106
rect 1935 1105 1939 1111
rect 1946 1109 1950 1113
rect 1954 1108 1958 1112
rect 1965 1110 1969 1116
rect 1984 1115 1988 1131
rect 1980 1108 1984 1112
rect 1932 1101 1942 1105
rect 1932 1094 1935 1096
rect 1939 1094 1942 1096
rect 1932 1093 1942 1094
rect 1950 1090 1954 1106
rect 1962 1102 1972 1103
rect 1962 1100 1965 1102
rect 1969 1100 1972 1102
rect 1962 1091 1972 1095
rect 1912 1083 1916 1087
rect 1920 1084 1924 1088
rect 1882 1064 1886 1081
rect 1894 1077 1904 1078
rect 1894 1075 1897 1077
rect 1901 1075 1904 1077
rect 1894 1066 1904 1070
rect 1886 1058 1890 1062
rect 1897 1060 1901 1066
rect 1916 1065 1920 1081
rect 1935 1080 1939 1086
rect 1946 1084 1950 1088
rect 1954 1083 1958 1087
rect 1965 1085 1969 1091
rect 1984 1090 1988 1106
rect 1980 1083 1984 1087
rect 1932 1076 1942 1080
rect 1932 1069 1935 1071
rect 1939 1069 1942 1071
rect 1932 1068 1942 1069
rect 1950 1065 1954 1081
rect 1962 1077 1972 1078
rect 1962 1075 1965 1077
rect 1969 1075 1972 1077
rect 1962 1066 1972 1070
rect 1912 1058 1916 1062
rect 1920 1059 1924 1063
rect 1882 1039 1886 1056
rect 1894 1052 1904 1053
rect 1894 1050 1897 1052
rect 1901 1050 1904 1052
rect 1894 1041 1904 1045
rect 1886 1033 1890 1037
rect 1897 1035 1901 1041
rect 1916 1040 1920 1056
rect 1935 1055 1939 1061
rect 1946 1059 1950 1063
rect 1954 1058 1958 1062
rect 1965 1060 1969 1066
rect 1984 1065 1988 1081
rect 1980 1058 1984 1062
rect 1932 1051 1942 1055
rect 1932 1044 1935 1046
rect 1939 1044 1942 1046
rect 1932 1043 1942 1044
rect 1950 1040 1954 1056
rect 1962 1052 1972 1053
rect 1962 1050 1965 1052
rect 1969 1050 1972 1052
rect 1962 1041 1972 1045
rect 1912 1033 1916 1037
rect 1920 1034 1924 1038
rect 938 1019 1865 1021
rect 1882 1019 1886 1031
rect 1894 1027 1904 1028
rect 1894 1025 1897 1027
rect 1901 1025 1904 1027
rect 938 1014 1886 1019
rect 1894 1016 1904 1020
rect 938 1006 1882 1014
rect 1886 1008 1890 1012
rect 1897 1010 1901 1016
rect 1916 1015 1920 1031
rect 1935 1030 1939 1036
rect 1946 1034 1950 1038
rect 1954 1033 1958 1037
rect 1965 1035 1969 1041
rect 1984 1040 1988 1056
rect 1980 1033 1984 1037
rect 1932 1026 1942 1030
rect 1932 1019 1935 1021
rect 1939 1019 1942 1021
rect 1932 1018 1942 1019
rect 1950 1015 1954 1031
rect 1962 1027 1972 1028
rect 1962 1025 1965 1027
rect 1969 1025 1972 1027
rect 1962 1016 1972 1020
rect 1912 1008 1916 1012
rect 1920 1009 1924 1013
rect 938 1005 1886 1006
rect 938 998 1865 1005
rect 910 997 1865 998
rect 909 993 1865 997
rect 1785 986 1865 993
rect -34 878 30 893
rect -34 670 4 878
rect 1828 785 1865 986
rect 1787 769 1865 785
rect 1795 745 1796 753
rect 1790 727 1804 733
rect -34 654 30 670
rect -34 524 4 654
rect 1828 555 1865 769
rect 1790 547 1865 555
rect -35 513 1790 524
rect -34 385 4 513
rect 1674 462 1702 466
rect 1745 459 1749 463
rect 1828 459 1865 547
rect 30 443 1865 459
rect -34 369 30 385
rect -34 237 4 369
rect 1828 311 1865 443
rect 1790 295 1865 311
rect 1790 267 1798 277
rect -34 220 30 237
rect -34 36 4 220
rect 1790 123 1817 131
rect 1828 110 1865 295
rect 1790 94 1865 110
rect -34 20 31 36
rect 1801 23 1807 25
rect 1780 12 1789 20
rect 1828 19 1865 94
rect 1882 989 1886 1005
rect 1894 1002 1904 1003
rect 1894 1000 1897 1002
rect 1901 1000 1904 1002
rect 1894 991 1904 995
rect 1886 983 1890 987
rect 1897 985 1901 991
rect 1916 990 1920 1006
rect 1935 1005 1939 1011
rect 1946 1009 1950 1013
rect 1954 1008 1958 1012
rect 1965 1010 1969 1016
rect 1984 1015 1988 1031
rect 1980 1008 1984 1012
rect 1932 1001 1942 1005
rect 1932 994 1935 996
rect 1939 994 1942 996
rect 1932 993 1942 994
rect 1950 990 1954 1006
rect 1962 1002 1972 1003
rect 1962 1000 1965 1002
rect 1969 1000 1972 1002
rect 1962 991 1972 995
rect 1912 983 1916 987
rect 1920 984 1924 988
rect 1882 964 1886 981
rect 1894 977 1904 978
rect 1894 975 1897 977
rect 1901 975 1904 977
rect 1894 966 1904 970
rect 1886 958 1890 962
rect 1897 960 1901 966
rect 1916 965 1920 981
rect 1935 980 1939 986
rect 1946 984 1950 988
rect 1954 983 1958 987
rect 1965 985 1969 991
rect 1984 990 1988 1006
rect 1980 983 1984 987
rect 1932 976 1942 980
rect 1932 969 1935 971
rect 1939 969 1942 971
rect 1932 968 1942 969
rect 1950 965 1954 981
rect 1962 977 1972 978
rect 1962 975 1965 977
rect 1969 975 1972 977
rect 1962 966 1972 970
rect 1912 958 1916 962
rect 1920 959 1924 963
rect 1882 939 1886 956
rect 1894 952 1904 953
rect 1894 950 1897 952
rect 1901 950 1904 952
rect 1894 941 1904 945
rect 1886 933 1890 937
rect 1897 935 1901 941
rect 1916 940 1920 956
rect 1935 955 1939 961
rect 1946 959 1950 963
rect 1954 958 1958 962
rect 1965 960 1969 966
rect 1984 965 1988 981
rect 1980 958 1984 962
rect 1932 951 1942 955
rect 1932 944 1935 946
rect 1939 944 1942 946
rect 1932 943 1942 944
rect 1950 940 1954 956
rect 1962 952 1972 953
rect 1962 950 1965 952
rect 1969 950 1972 952
rect 1962 941 1972 945
rect 1912 933 1916 937
rect 1920 934 1924 938
rect 1882 914 1886 931
rect 1894 927 1904 928
rect 1894 925 1897 927
rect 1901 925 1904 927
rect 1894 916 1904 920
rect 1886 908 1890 912
rect 1897 910 1901 916
rect 1916 915 1920 931
rect 1935 930 1939 936
rect 1946 934 1950 938
rect 1954 933 1958 937
rect 1965 935 1969 941
rect 1984 940 1988 956
rect 1980 933 1984 937
rect 1932 926 1942 930
rect 1932 919 1935 921
rect 1939 919 1942 921
rect 1932 918 1942 919
rect 1950 915 1954 931
rect 1962 927 1972 928
rect 1962 925 1965 927
rect 1969 925 1972 927
rect 1962 916 1972 920
rect 1912 908 1916 912
rect 1920 909 1924 913
rect 1882 889 1886 906
rect 1894 902 1904 903
rect 1894 900 1897 902
rect 1901 900 1904 902
rect 1894 891 1904 895
rect 1886 883 1890 887
rect 1897 885 1901 891
rect 1916 890 1920 906
rect 1935 905 1939 911
rect 1946 909 1950 913
rect 1954 908 1958 912
rect 1965 910 1969 916
rect 1984 915 1988 931
rect 1980 908 1984 912
rect 1932 901 1942 905
rect 1932 894 1935 896
rect 1939 894 1942 896
rect 1932 893 1942 894
rect 1950 890 1954 906
rect 1962 902 1972 903
rect 1962 900 1965 902
rect 1969 900 1972 902
rect 1962 891 1972 895
rect 1912 883 1916 887
rect 1920 884 1924 888
rect 1882 864 1886 881
rect 1894 877 1904 878
rect 1894 875 1897 877
rect 1901 875 1904 877
rect 1894 866 1904 870
rect 1886 858 1890 862
rect 1897 860 1901 866
rect 1916 865 1920 881
rect 1935 880 1939 886
rect 1946 884 1950 888
rect 1954 883 1958 887
rect 1965 885 1969 891
rect 1984 890 1988 906
rect 1980 883 1984 887
rect 1932 876 1942 880
rect 1932 869 1935 871
rect 1939 869 1942 871
rect 1932 868 1942 869
rect 1950 865 1954 881
rect 1962 877 1972 878
rect 1962 875 1965 877
rect 1969 875 1972 877
rect 1962 866 1972 870
rect 1912 858 1916 862
rect 1920 859 1924 863
rect 1882 839 1886 856
rect 1894 852 1904 853
rect 1894 850 1897 852
rect 1901 850 1904 852
rect 1894 841 1904 845
rect 1886 833 1890 837
rect 1897 835 1901 841
rect 1916 840 1920 856
rect 1935 855 1939 861
rect 1946 859 1950 863
rect 1954 858 1958 862
rect 1965 860 1969 866
rect 1984 865 1988 881
rect 1980 858 1984 862
rect 1932 851 1942 855
rect 1932 844 1935 846
rect 1939 844 1942 846
rect 1932 843 1942 844
rect 1950 840 1954 856
rect 1962 852 1972 853
rect 1962 850 1965 852
rect 1969 850 1972 852
rect 1962 841 1972 845
rect 1912 833 1916 837
rect 1920 834 1924 838
rect 1882 814 1886 831
rect 1894 827 1904 828
rect 1894 825 1897 827
rect 1901 825 1904 827
rect 1894 816 1904 820
rect 1886 808 1890 812
rect 1897 810 1901 816
rect 1916 815 1920 831
rect 1935 830 1939 836
rect 1946 834 1950 838
rect 1954 833 1958 837
rect 1965 835 1969 841
rect 1984 840 1988 856
rect 1980 833 1984 837
rect 1932 826 1942 830
rect 1932 819 1935 821
rect 1939 819 1942 821
rect 1932 818 1942 819
rect 1950 815 1954 831
rect 1962 827 1972 828
rect 1962 825 1965 827
rect 1969 825 1972 827
rect 1962 816 1972 820
rect 1912 808 1916 812
rect 1920 809 1924 813
rect 1882 789 1886 806
rect 1894 802 1904 803
rect 1894 800 1897 802
rect 1901 800 1904 802
rect 1894 791 1904 795
rect 1886 783 1890 787
rect 1897 785 1901 791
rect 1916 790 1920 806
rect 1935 805 1939 811
rect 1946 809 1950 813
rect 1954 808 1958 812
rect 1965 810 1969 816
rect 1984 815 1988 831
rect 1980 808 1984 812
rect 1932 801 1942 805
rect 1932 794 1935 796
rect 1939 794 1942 796
rect 1932 793 1942 794
rect 1950 790 1954 806
rect 1962 802 1972 803
rect 1962 800 1965 802
rect 1969 800 1972 802
rect 1962 791 1972 795
rect 1912 783 1916 787
rect 1920 784 1924 788
rect 1882 764 1886 781
rect 1894 777 1904 778
rect 1894 775 1897 777
rect 1901 775 1904 777
rect 1894 766 1904 770
rect 1886 758 1890 762
rect 1897 760 1901 766
rect 1916 765 1920 781
rect 1935 780 1939 786
rect 1946 784 1950 788
rect 1954 783 1958 787
rect 1965 785 1969 791
rect 1984 790 1988 806
rect 1980 783 1984 787
rect 1932 776 1942 780
rect 1932 769 1935 771
rect 1939 769 1942 771
rect 1932 768 1942 769
rect 1950 765 1954 781
rect 1962 777 1972 778
rect 1962 775 1965 777
rect 1969 775 1972 777
rect 1962 766 1972 770
rect 1912 758 1916 762
rect 1920 759 1924 763
rect 1882 739 1886 756
rect 1894 752 1904 753
rect 1894 750 1897 752
rect 1901 750 1904 752
rect 1894 741 1904 745
rect 1886 733 1890 737
rect 1897 735 1901 741
rect 1916 740 1920 756
rect 1935 755 1939 761
rect 1946 759 1950 763
rect 1954 758 1958 762
rect 1965 760 1969 766
rect 1984 765 1988 781
rect 1980 758 1984 762
rect 1932 751 1942 755
rect 1932 744 1935 746
rect 1939 744 1942 746
rect 1932 743 1942 744
rect 1950 740 1954 756
rect 1962 752 1972 753
rect 1962 750 1965 752
rect 1969 750 1972 752
rect 1962 741 1972 745
rect 1912 733 1916 737
rect 1920 734 1924 738
rect 1882 714 1886 731
rect 1894 727 1904 728
rect 1894 725 1897 727
rect 1901 725 1904 727
rect 1894 716 1904 720
rect 1886 708 1890 712
rect 1897 710 1901 716
rect 1916 715 1920 731
rect 1935 730 1939 736
rect 1946 734 1950 738
rect 1954 733 1958 737
rect 1965 735 1969 741
rect 1984 740 1988 756
rect 1980 733 1984 737
rect 1932 726 1942 730
rect 1932 719 1935 721
rect 1939 719 1942 721
rect 1932 718 1942 719
rect 1950 715 1954 731
rect 1962 727 1972 728
rect 1962 725 1965 727
rect 1969 725 1972 727
rect 1962 716 1972 720
rect 1912 708 1916 712
rect 1920 709 1924 713
rect 1882 689 1886 706
rect 1894 702 1904 703
rect 1894 700 1897 702
rect 1901 700 1904 702
rect 1894 691 1904 695
rect 1886 683 1890 687
rect 1897 685 1901 691
rect 1916 690 1920 706
rect 1935 705 1939 711
rect 1946 709 1950 713
rect 1954 708 1958 712
rect 1965 710 1969 716
rect 1984 715 1988 731
rect 1980 708 1984 712
rect 1932 701 1942 705
rect 1932 694 1935 696
rect 1939 694 1942 696
rect 1932 693 1942 694
rect 1950 690 1954 706
rect 1962 702 1972 703
rect 1962 700 1965 702
rect 1969 700 1972 702
rect 1962 691 1972 695
rect 1912 683 1916 687
rect 1920 684 1924 688
rect 1882 664 1886 681
rect 1894 677 1904 678
rect 1894 675 1897 677
rect 1901 675 1904 677
rect 1894 666 1904 670
rect 1886 658 1890 662
rect 1897 660 1901 666
rect 1916 665 1920 681
rect 1935 680 1939 686
rect 1946 684 1950 688
rect 1954 683 1958 687
rect 1965 685 1969 691
rect 1984 690 1988 706
rect 1980 683 1984 687
rect 1932 676 1942 680
rect 1932 669 1935 671
rect 1939 669 1942 671
rect 1932 668 1942 669
rect 1950 665 1954 681
rect 1962 677 1972 678
rect 1962 675 1965 677
rect 1969 675 1972 677
rect 1962 666 1972 670
rect 1912 658 1916 662
rect 1920 659 1924 663
rect 1882 639 1886 656
rect 1894 652 1904 653
rect 1894 650 1897 652
rect 1901 650 1904 652
rect 1894 641 1904 645
rect 1886 633 1890 637
rect 1897 635 1901 641
rect 1916 640 1920 656
rect 1935 655 1939 661
rect 1946 659 1950 663
rect 1954 658 1958 662
rect 1965 660 1969 666
rect 1984 665 1988 681
rect 1980 658 1984 662
rect 1932 651 1942 655
rect 1932 644 1935 646
rect 1939 644 1942 646
rect 1932 643 1942 644
rect 1950 640 1954 656
rect 1962 652 1972 653
rect 1962 650 1965 652
rect 1969 650 1972 652
rect 1962 641 1972 645
rect 1912 633 1916 637
rect 1920 634 1924 638
rect 1882 614 1886 631
rect 1894 627 1904 628
rect 1894 625 1897 627
rect 1901 625 1904 627
rect 1894 616 1904 620
rect 1886 608 1890 612
rect 1897 610 1901 616
rect 1916 615 1920 631
rect 1935 630 1939 636
rect 1946 634 1950 638
rect 1954 633 1958 637
rect 1965 635 1969 641
rect 1984 640 1988 656
rect 1980 633 1984 637
rect 1932 626 1942 630
rect 1932 619 1935 621
rect 1939 619 1942 621
rect 1932 618 1942 619
rect 1950 615 1954 631
rect 1962 627 1972 628
rect 1962 625 1965 627
rect 1969 625 1972 627
rect 1962 616 1972 620
rect 1912 608 1916 612
rect 1920 609 1924 613
rect 1882 589 1886 606
rect 1894 602 1904 603
rect 1894 600 1897 602
rect 1901 600 1904 602
rect 1894 591 1904 595
rect 1886 583 1890 587
rect 1897 585 1901 591
rect 1916 590 1920 606
rect 1935 605 1939 611
rect 1946 609 1950 613
rect 1954 608 1958 612
rect 1965 610 1969 616
rect 1984 615 1988 631
rect 1980 608 1984 612
rect 1932 601 1942 605
rect 1932 594 1935 596
rect 1939 594 1942 596
rect 1932 593 1942 594
rect 1950 590 1954 606
rect 1962 602 1972 603
rect 1962 600 1965 602
rect 1969 600 1972 602
rect 1962 591 1972 595
rect 1912 583 1916 587
rect 1920 584 1924 588
rect 1882 564 1886 581
rect 1894 577 1904 578
rect 1894 575 1897 577
rect 1901 575 1904 577
rect 1894 566 1904 570
rect 1886 558 1890 562
rect 1897 560 1901 566
rect 1916 565 1920 581
rect 1935 580 1939 586
rect 1946 584 1950 588
rect 1954 583 1958 587
rect 1965 585 1969 591
rect 1984 590 1988 606
rect 1980 583 1984 587
rect 1932 576 1942 580
rect 1932 569 1935 571
rect 1939 569 1942 571
rect 1932 568 1942 569
rect 1950 565 1954 581
rect 1962 577 1972 578
rect 1962 575 1965 577
rect 1969 575 1972 577
rect 1962 566 1972 570
rect 1912 558 1916 562
rect 1920 559 1924 563
rect 1882 539 1886 556
rect 1894 552 1904 553
rect 1894 550 1897 552
rect 1901 550 1904 552
rect 1894 541 1904 545
rect 1886 533 1890 537
rect 1897 535 1901 541
rect 1916 540 1920 556
rect 1935 555 1939 561
rect 1946 559 1950 563
rect 1954 558 1958 562
rect 1965 560 1969 566
rect 1984 565 1988 581
rect 1980 558 1984 562
rect 1932 551 1942 555
rect 1932 544 1935 546
rect 1939 544 1942 546
rect 1932 543 1942 544
rect 1950 540 1954 556
rect 1962 552 1972 553
rect 1962 550 1965 552
rect 1969 550 1972 552
rect 1962 541 1972 545
rect 1912 533 1916 537
rect 1920 534 1924 538
rect 1882 514 1886 531
rect 1894 527 1904 528
rect 1894 525 1897 527
rect 1901 525 1904 527
rect 1894 516 1904 520
rect 1886 508 1890 512
rect 1897 510 1901 516
rect 1916 515 1920 531
rect 1935 530 1939 536
rect 1946 534 1950 538
rect 1954 533 1958 537
rect 1965 535 1969 541
rect 1984 540 1988 556
rect 1980 533 1984 537
rect 1932 526 1942 530
rect 1932 519 1935 521
rect 1939 519 1942 521
rect 1932 518 1942 519
rect 1950 515 1954 531
rect 1962 527 1972 528
rect 1962 525 1965 527
rect 1969 525 1972 527
rect 1962 516 1972 520
rect 1912 508 1916 512
rect 1920 509 1924 513
rect 1882 489 1886 506
rect 1894 502 1904 503
rect 1894 500 1897 502
rect 1901 500 1904 502
rect 1894 491 1904 495
rect 1886 483 1890 487
rect 1897 485 1901 491
rect 1916 490 1920 506
rect 1935 505 1939 511
rect 1946 509 1950 513
rect 1954 508 1958 512
rect 1965 510 1969 516
rect 1984 515 1988 531
rect 1980 508 1984 512
rect 1932 501 1942 505
rect 1932 494 1935 496
rect 1939 494 1942 496
rect 1932 493 1942 494
rect 1950 490 1954 506
rect 1962 502 1972 503
rect 1962 500 1965 502
rect 1969 500 1972 502
rect 1962 491 1972 495
rect 1912 483 1916 487
rect 1920 484 1924 488
rect 1882 464 1886 481
rect 1894 477 1904 478
rect 1894 475 1897 477
rect 1901 475 1904 477
rect 1894 466 1904 470
rect 1886 458 1890 462
rect 1897 460 1901 466
rect 1916 465 1920 481
rect 1935 480 1939 486
rect 1946 484 1950 488
rect 1954 483 1958 487
rect 1965 485 1969 491
rect 1984 490 1988 506
rect 1980 483 1984 487
rect 1932 476 1942 480
rect 1932 469 1935 471
rect 1939 469 1942 471
rect 1932 468 1942 469
rect 1950 465 1954 481
rect 1962 477 1972 478
rect 1962 475 1965 477
rect 1969 475 1972 477
rect 1962 466 1972 470
rect 1912 458 1916 462
rect 1920 459 1924 463
rect 1882 439 1886 456
rect 1894 452 1904 453
rect 1894 450 1897 452
rect 1901 450 1904 452
rect 1894 441 1904 445
rect 1886 433 1890 437
rect 1897 435 1901 441
rect 1916 440 1920 456
rect 1935 455 1939 461
rect 1946 459 1950 463
rect 1954 458 1958 462
rect 1965 460 1969 466
rect 1984 465 1988 481
rect 1980 458 1984 462
rect 1932 451 1942 455
rect 1932 444 1935 446
rect 1939 444 1942 446
rect 1932 443 1942 444
rect 1950 440 1954 456
rect 1962 452 1972 453
rect 1962 450 1965 452
rect 1969 450 1972 452
rect 1962 441 1972 445
rect 1912 433 1916 437
rect 1920 434 1924 438
rect 1882 414 1886 431
rect 1894 427 1904 428
rect 1894 425 1897 427
rect 1901 425 1904 427
rect 1894 416 1904 420
rect 1886 408 1890 412
rect 1897 410 1901 416
rect 1916 415 1920 431
rect 1935 430 1939 436
rect 1946 434 1950 438
rect 1954 433 1958 437
rect 1965 435 1969 441
rect 1984 440 1988 456
rect 1980 433 1984 437
rect 1932 426 1942 430
rect 1932 419 1935 421
rect 1939 419 1942 421
rect 1932 418 1942 419
rect 1950 415 1954 431
rect 1962 427 1972 428
rect 1962 425 1965 427
rect 1969 425 1972 427
rect 1962 416 1972 420
rect 1912 408 1916 412
rect 1920 409 1924 413
rect 1882 389 1886 406
rect 1894 402 1904 403
rect 1894 400 1897 402
rect 1901 400 1904 402
rect 1894 391 1904 395
rect 1886 383 1890 387
rect 1897 385 1901 391
rect 1916 390 1920 406
rect 1935 405 1939 411
rect 1946 409 1950 413
rect 1954 408 1958 412
rect 1965 410 1969 416
rect 1984 415 1988 431
rect 1980 408 1984 412
rect 1932 401 1942 405
rect 1932 394 1935 396
rect 1939 394 1942 396
rect 1932 393 1942 394
rect 1950 390 1954 406
rect 1962 402 1972 403
rect 1962 400 1965 402
rect 1969 400 1972 402
rect 1962 391 1972 395
rect 1912 383 1916 387
rect 1920 384 1924 388
rect 1882 364 1886 381
rect 1894 377 1904 378
rect 1894 375 1897 377
rect 1901 375 1904 377
rect 1894 366 1904 370
rect 1886 358 1890 362
rect 1897 360 1901 366
rect 1916 365 1920 381
rect 1935 380 1939 386
rect 1946 384 1950 388
rect 1954 383 1958 387
rect 1965 385 1969 391
rect 1984 390 1988 406
rect 1980 383 1984 387
rect 1932 376 1942 380
rect 1932 369 1935 371
rect 1939 369 1942 371
rect 1932 368 1942 369
rect 1950 365 1954 381
rect 1962 377 1972 378
rect 1962 375 1965 377
rect 1969 375 1972 377
rect 1962 366 1972 370
rect 1912 358 1916 362
rect 1920 359 1924 363
rect 1882 339 1886 356
rect 1894 352 1904 353
rect 1894 350 1897 352
rect 1901 350 1904 352
rect 1894 341 1904 345
rect 1886 333 1890 337
rect 1897 335 1901 341
rect 1916 340 1920 356
rect 1935 355 1939 361
rect 1946 359 1950 363
rect 1954 358 1958 362
rect 1965 360 1969 366
rect 1984 365 1988 381
rect 1980 358 1984 362
rect 1932 351 1942 355
rect 1932 344 1935 346
rect 1939 344 1942 346
rect 1932 343 1942 344
rect 1950 340 1954 356
rect 1962 352 1972 353
rect 1962 350 1965 352
rect 1969 350 1972 352
rect 1962 341 1972 345
rect 1912 333 1916 337
rect 1920 334 1924 338
rect 1882 314 1886 331
rect 1894 327 1904 328
rect 1894 325 1897 327
rect 1901 325 1904 327
rect 1894 316 1904 320
rect 1886 308 1890 312
rect 1897 310 1901 316
rect 1916 315 1920 331
rect 1935 330 1939 336
rect 1946 334 1950 338
rect 1954 333 1958 337
rect 1965 335 1969 341
rect 1984 340 1988 356
rect 1980 333 1984 337
rect 1932 326 1942 330
rect 1932 319 1935 321
rect 1939 319 1942 321
rect 1932 318 1942 319
rect 1950 315 1954 331
rect 1962 327 1972 328
rect 1962 325 1965 327
rect 1969 325 1972 327
rect 1962 316 1972 320
rect 1912 308 1916 312
rect 1920 309 1924 313
rect 1882 289 1886 306
rect 1894 302 1904 303
rect 1894 300 1897 302
rect 1901 300 1904 302
rect 1894 291 1904 295
rect 1886 283 1890 287
rect 1897 285 1901 291
rect 1916 290 1920 306
rect 1935 305 1939 311
rect 1946 309 1950 313
rect 1954 308 1958 312
rect 1965 310 1969 316
rect 1984 315 1988 331
rect 1980 308 1984 312
rect 1932 301 1942 305
rect 1932 294 1935 296
rect 1939 294 1942 296
rect 1932 293 1942 294
rect 1950 290 1954 306
rect 1962 302 1972 303
rect 1962 300 1965 302
rect 1969 300 1972 302
rect 1962 291 1972 295
rect 1912 283 1916 287
rect 1920 284 1924 288
rect 1882 264 1886 281
rect 1894 277 1904 278
rect 1894 275 1897 277
rect 1901 275 1904 277
rect 1894 266 1904 270
rect 1886 258 1890 262
rect 1897 260 1901 266
rect 1916 265 1920 281
rect 1935 280 1939 286
rect 1946 284 1950 288
rect 1954 283 1958 287
rect 1965 285 1969 291
rect 1984 290 1988 306
rect 1980 283 1984 287
rect 1932 276 1942 280
rect 1932 269 1935 271
rect 1939 269 1942 271
rect 1932 268 1942 269
rect 1950 265 1954 281
rect 1962 277 1972 278
rect 1962 275 1965 277
rect 1969 275 1972 277
rect 1962 266 1972 270
rect 1912 258 1916 262
rect 1920 259 1924 263
rect 1882 239 1886 256
rect 1894 252 1904 253
rect 1894 250 1897 252
rect 1901 250 1904 252
rect 1894 241 1904 245
rect 1886 233 1890 237
rect 1897 235 1901 241
rect 1916 240 1920 256
rect 1935 255 1939 261
rect 1946 259 1950 263
rect 1954 258 1958 262
rect 1965 260 1969 266
rect 1984 265 1988 281
rect 1980 258 1984 262
rect 1932 251 1942 255
rect 1932 244 1935 246
rect 1939 244 1942 246
rect 1932 243 1942 244
rect 1950 240 1954 256
rect 1962 252 1972 253
rect 1962 250 1965 252
rect 1969 250 1972 252
rect 1962 241 1972 245
rect 1912 233 1916 237
rect 1920 234 1924 238
rect 1882 214 1886 231
rect 1894 227 1904 228
rect 1894 225 1897 227
rect 1901 225 1904 227
rect 1894 216 1904 220
rect 1886 208 1890 212
rect 1897 210 1901 216
rect 1916 215 1920 231
rect 1935 230 1939 236
rect 1946 234 1950 238
rect 1954 233 1958 237
rect 1965 235 1969 241
rect 1984 240 1988 256
rect 1980 233 1984 237
rect 1932 226 1942 230
rect 1932 219 1935 221
rect 1939 219 1942 221
rect 1932 218 1942 219
rect 1950 215 1954 231
rect 1962 227 1972 228
rect 1962 225 1965 227
rect 1969 225 1972 227
rect 1962 216 1972 220
rect 1912 208 1916 212
rect 1920 209 1924 213
rect 1882 189 1886 206
rect 1894 202 1904 203
rect 1894 200 1897 202
rect 1901 200 1904 202
rect 1894 191 1904 195
rect 1886 183 1890 187
rect 1897 185 1901 191
rect 1916 190 1920 206
rect 1935 205 1939 211
rect 1946 209 1950 213
rect 1954 208 1958 212
rect 1965 210 1969 216
rect 1984 215 1988 231
rect 1980 208 1984 212
rect 1932 201 1942 205
rect 1932 194 1935 196
rect 1939 194 1942 196
rect 1932 193 1942 194
rect 1950 190 1954 206
rect 1962 202 1972 203
rect 1962 200 1965 202
rect 1969 200 1972 202
rect 1962 191 1972 195
rect 1912 183 1916 187
rect 1920 184 1924 188
rect 1882 164 1886 181
rect 1894 177 1904 178
rect 1894 175 1897 177
rect 1901 175 1904 177
rect 1894 166 1904 170
rect 1886 158 1890 162
rect 1897 160 1901 166
rect 1916 165 1920 181
rect 1935 180 1939 186
rect 1946 184 1950 188
rect 1954 183 1958 187
rect 1965 185 1969 191
rect 1984 190 1988 206
rect 1980 183 1984 187
rect 1932 176 1942 180
rect 1932 169 1935 171
rect 1939 169 1942 171
rect 1932 168 1942 169
rect 1950 165 1954 181
rect 1962 177 1972 178
rect 1962 175 1965 177
rect 1969 175 1972 177
rect 1962 166 1972 170
rect 1912 158 1916 162
rect 1920 159 1924 163
rect 1882 139 1886 156
rect 1894 152 1904 153
rect 1894 150 1897 152
rect 1901 150 1904 152
rect 1894 141 1904 145
rect 1886 133 1890 137
rect 1897 135 1901 141
rect 1916 140 1920 156
rect 1935 155 1939 161
rect 1946 159 1950 163
rect 1954 158 1958 162
rect 1965 160 1969 166
rect 1984 165 1988 181
rect 1980 158 1984 162
rect 1932 151 1942 155
rect 1932 144 1935 146
rect 1939 144 1942 146
rect 1932 143 1942 144
rect 1950 140 1954 156
rect 1962 152 1972 153
rect 1962 150 1965 152
rect 1969 150 1972 152
rect 1962 141 1972 145
rect 1912 133 1916 137
rect 1920 134 1924 138
rect 1882 114 1886 131
rect 1894 127 1904 128
rect 1894 125 1897 127
rect 1901 125 1904 127
rect 1894 116 1904 120
rect 1886 108 1890 112
rect 1897 110 1901 116
rect 1916 115 1920 131
rect 1935 130 1939 136
rect 1946 134 1950 138
rect 1954 133 1958 137
rect 1965 135 1969 141
rect 1984 140 1988 156
rect 1980 133 1984 137
rect 1932 126 1942 130
rect 1932 119 1935 121
rect 1939 119 1942 121
rect 1932 118 1942 119
rect 1950 115 1954 131
rect 1962 127 1972 128
rect 1962 125 1965 127
rect 1969 125 1972 127
rect 1962 116 1972 120
rect 1912 108 1916 112
rect 1920 109 1924 113
rect 1882 89 1886 106
rect 1894 102 1904 103
rect 1894 100 1897 102
rect 1901 100 1904 102
rect 1894 91 1904 95
rect 1886 83 1890 87
rect 1897 85 1901 91
rect 1916 90 1920 106
rect 1935 105 1939 111
rect 1946 109 1950 113
rect 1954 108 1958 112
rect 1965 110 1969 116
rect 1984 115 1988 131
rect 1980 108 1984 112
rect 1932 101 1942 105
rect 1932 94 1935 96
rect 1939 94 1942 96
rect 1932 93 1942 94
rect 1950 90 1954 106
rect 1962 102 1972 103
rect 1962 100 1965 102
rect 1969 100 1972 102
rect 1962 91 1972 95
rect 1912 83 1916 87
rect 1920 84 1924 88
rect 1882 64 1886 81
rect 1894 77 1904 78
rect 1894 75 1897 77
rect 1901 75 1904 77
rect 1894 66 1904 70
rect 1886 58 1890 62
rect 1897 60 1901 66
rect 1916 65 1920 81
rect 1935 80 1939 86
rect 1946 84 1950 88
rect 1954 83 1958 87
rect 1965 85 1969 91
rect 1984 90 1988 106
rect 1980 83 1984 87
rect 1932 76 1942 80
rect 1932 69 1935 71
rect 1939 69 1942 71
rect 1932 68 1942 69
rect 1950 65 1954 81
rect 1962 77 1972 78
rect 1962 75 1965 77
rect 1969 75 1972 77
rect 1962 66 1972 70
rect 1912 58 1916 62
rect 1920 59 1924 63
rect 1882 39 1886 56
rect 1894 52 1904 53
rect 1894 50 1897 52
rect 1901 50 1904 52
rect 1894 41 1904 45
rect 1886 33 1890 37
rect 1897 35 1901 41
rect 1916 40 1920 56
rect 1935 55 1939 61
rect 1946 59 1950 63
rect 1954 58 1958 62
rect 1965 60 1969 66
rect 1984 65 1988 81
rect 1980 58 1984 62
rect 1932 51 1942 55
rect 1932 44 1935 46
rect 1939 44 1942 46
rect 1932 43 1942 44
rect 1950 40 1954 56
rect 1962 52 1972 53
rect 1962 50 1965 52
rect 1969 50 1972 52
rect 1962 41 1972 45
rect 1912 33 1916 37
rect 1920 34 1924 38
rect 1882 23 1886 31
rect 1894 27 1904 28
rect 1894 25 1897 27
rect 1901 25 1904 27
rect 1916 20 1920 31
rect 1935 30 1939 36
rect 1946 34 1950 38
rect 1954 33 1958 37
rect 1965 35 1969 41
rect 1984 40 1988 56
rect 1980 33 1984 37
rect 1932 26 1942 30
rect 1950 23 1954 31
rect 1962 27 1972 28
rect 1962 25 1965 27
rect 1969 25 1972 27
rect 1984 20 1988 31
rect 1916 15 1988 20
rect 1933 12 1943 15
rect 1780 3 1947 12
<< metal2 >>
rect 12 1039 20 1880
rect 43 1833 49 1864
rect 43 1823 49 1828
rect 153 1834 159 1864
rect 153 1823 159 1829
rect 263 1833 269 1864
rect 263 1823 269 1828
rect 373 1834 379 1864
rect 373 1823 379 1829
rect 483 1834 489 1864
rect 483 1823 489 1829
rect 593 1833 599 1864
rect 593 1823 599 1828
rect 703 1833 709 1864
rect 703 1823 709 1828
rect 813 1833 819 1864
rect 813 1823 819 1828
rect 920 1643 928 2006
rect 1011 2013 1110 2017
rect 1011 1953 1024 2013
rect 925 1635 928 1643
rect 917 1336 925 1617
rect 1104 1605 1110 2013
rect 1121 2012 1220 2017
rect 1121 1956 1134 2012
rect 1214 1605 1220 2012
rect 1231 2012 1330 2017
rect 1231 1956 1244 2012
rect 1324 1605 1330 2012
rect 1341 2012 1440 2017
rect 1341 1956 1354 2012
rect 1104 1599 1124 1605
rect 1214 1599 1229 1605
rect 1324 1599 1344 1605
rect 995 1565 1011 1571
rect 935 1446 991 1454
rect 917 1328 949 1336
rect 910 1316 933 1320
rect 925 1036 933 1316
rect 941 1052 949 1328
rect 981 1226 991 1446
rect 995 1167 1001 1565
rect 1010 1544 1111 1550
rect 1118 1544 1222 1548
rect 1105 1168 1111 1544
rect 1216 1168 1222 1544
rect 1229 1542 1333 1548
rect 1327 1169 1333 1542
rect 1424 1381 1430 1657
rect 1434 1605 1440 2012
rect 1451 2012 1550 2017
rect 1451 1956 1464 2012
rect 1544 1605 1550 2012
rect 1561 1956 1574 2017
rect 1662 1889 1696 1897
rect 1661 1743 1682 1753
rect 1434 1599 1454 1605
rect 1544 1599 1564 1605
rect 1546 1333 1554 1463
rect 1674 1411 1682 1743
rect 1686 1348 1696 1889
rect 1657 1324 1673 1332
rect 1658 1316 1673 1324
rect 1786 1264 1804 1268
rect 1778 1256 1796 1260
rect 1778 1158 1812 1162
rect 1755 1135 1865 1139
rect 1754 1105 1828 1112
rect 1779 1097 1789 1101
rect 1005 1088 1869 1092
rect 941 1044 979 1052
rect 925 1028 979 1036
rect 1005 994 1011 1088
rect 1115 1080 1869 1084
rect 1115 994 1121 1080
rect 1225 1072 1869 1076
rect 1225 994 1231 1072
rect 1335 1064 1869 1068
rect 1335 994 1341 1064
rect 1445 1056 1869 1060
rect 1445 994 1451 1056
rect 1555 1048 1869 1052
rect 1555 994 1561 1048
rect 1665 1040 1869 1044
rect 1665 994 1671 1040
rect 1752 1028 1762 1036
rect 1774 1032 1869 1036
rect 1774 994 1780 1032
rect 1796 753 1800 1024
rect 1804 733 1808 1024
rect 1812 501 1816 1024
rect 1790 493 1812 501
rect 1820 469 1824 1024
rect 1790 466 1820 469
rect 1717 457 1721 465
rect 1794 462 1820 466
rect 1695 452 1721 457
rect 1695 432 1701 452
rect 1828 277 1836 1024
rect 1806 267 1812 277
rect 1820 267 1836 277
rect 1801 31 1807 267
rect 1844 131 1852 1024
rect 1823 123 1852 131
rect 81 17 94 20
rect 81 -21 94 11
rect 191 17 204 20
rect 191 -21 204 11
rect 301 17 314 20
rect 301 -21 314 11
rect 411 17 424 20
rect 411 -21 424 11
rect 521 17 534 20
rect 521 -21 534 11
rect 631 17 644 20
rect 631 -21 644 11
rect 741 17 754 20
rect 741 -21 754 11
rect 851 17 864 20
rect 851 -21 864 11
rect 961 17 974 20
rect 961 -21 974 11
rect 1071 17 1084 20
rect 1071 -21 1084 11
rect 1181 17 1194 20
rect 1181 -21 1194 11
rect 1291 17 1304 20
rect 1291 -21 1304 11
rect 1401 17 1414 20
rect 1401 -21 1414 11
rect 1511 17 1524 20
rect 1511 -21 1524 11
rect 1621 17 1634 20
rect 1621 -21 1634 11
rect 1731 17 1744 20
rect 1731 -21 1744 11
<< ntransistor >>
rect 1890 2013 1894 2015
rect 1890 2005 1894 2007
rect 1942 2014 1946 2016
rect 1942 2006 1946 2008
rect 1958 2013 1962 2015
rect 1958 2005 1962 2007
rect 1890 1988 1894 1990
rect 1890 1980 1894 1982
rect 1942 1989 1946 1991
rect 1942 1981 1946 1983
rect 1958 1988 1962 1990
rect 1958 1980 1962 1982
rect 1890 1963 1894 1965
rect 1890 1955 1894 1957
rect 1942 1964 1946 1966
rect 1942 1956 1946 1958
rect 1958 1963 1962 1965
rect 1958 1955 1962 1957
rect 1890 1938 1894 1940
rect 1890 1930 1894 1932
rect 1942 1939 1946 1941
rect 1942 1931 1946 1933
rect 1958 1938 1962 1940
rect 1958 1930 1962 1932
rect 1890 1913 1894 1915
rect 1890 1905 1894 1907
rect 1942 1914 1946 1916
rect 1942 1906 1946 1908
rect 1958 1913 1962 1915
rect 1958 1905 1962 1907
rect 1890 1888 1894 1890
rect 1890 1880 1894 1882
rect 1942 1889 1946 1891
rect 1942 1881 1946 1883
rect 1958 1888 1962 1890
rect 1958 1880 1962 1882
rect 1890 1863 1894 1865
rect 1890 1855 1894 1857
rect 1942 1864 1946 1866
rect 1942 1856 1946 1858
rect 1958 1863 1962 1865
rect 1958 1855 1962 1857
rect 1890 1838 1894 1840
rect 1890 1830 1894 1832
rect 1942 1839 1946 1841
rect 1942 1831 1946 1833
rect 1958 1838 1962 1840
rect 1958 1830 1962 1832
rect 1890 1813 1894 1815
rect 1890 1805 1894 1807
rect 1942 1814 1946 1816
rect 1942 1806 1946 1808
rect 1958 1813 1962 1815
rect 1958 1805 1962 1807
rect 1890 1788 1894 1790
rect 1890 1780 1894 1782
rect 1942 1789 1946 1791
rect 1942 1781 1946 1783
rect 1958 1788 1962 1790
rect 1958 1780 1962 1782
rect 1890 1763 1894 1765
rect 1890 1755 1894 1757
rect 1942 1764 1946 1766
rect 1942 1756 1946 1758
rect 1958 1763 1962 1765
rect 1958 1755 1962 1757
rect 1890 1738 1894 1740
rect 1890 1730 1894 1732
rect 1942 1739 1946 1741
rect 1942 1731 1946 1733
rect 1958 1738 1962 1740
rect 1958 1730 1962 1732
rect 1890 1713 1894 1715
rect 1890 1705 1894 1707
rect 1942 1714 1946 1716
rect 1942 1706 1946 1708
rect 1958 1713 1962 1715
rect 1958 1705 1962 1707
rect 1890 1688 1894 1690
rect 1890 1680 1894 1682
rect 1942 1689 1946 1691
rect 1942 1681 1946 1683
rect 1958 1688 1962 1690
rect 1958 1680 1962 1682
rect 1890 1663 1894 1665
rect 1890 1655 1894 1657
rect 1942 1664 1946 1666
rect 1942 1656 1946 1658
rect 1958 1663 1962 1665
rect 1958 1655 1962 1657
rect 1890 1638 1894 1640
rect 1890 1630 1894 1632
rect 1942 1639 1946 1641
rect 1942 1631 1946 1633
rect 1958 1638 1962 1640
rect 1958 1630 1962 1632
rect 1890 1613 1894 1615
rect 1890 1605 1894 1607
rect 1942 1614 1946 1616
rect 1942 1606 1946 1608
rect 1958 1613 1962 1615
rect 1958 1605 1962 1607
rect 1890 1588 1894 1590
rect 1890 1580 1894 1582
rect 1942 1589 1946 1591
rect 1942 1581 1946 1583
rect 1958 1588 1962 1590
rect 1958 1580 1962 1582
rect 1890 1563 1894 1565
rect 1890 1555 1894 1557
rect 1942 1564 1946 1566
rect 1942 1556 1946 1558
rect 1958 1563 1962 1565
rect 1958 1555 1962 1557
rect 1890 1538 1894 1540
rect 1890 1530 1894 1532
rect 1942 1539 1946 1541
rect 1942 1531 1946 1533
rect 1958 1538 1962 1540
rect 1958 1530 1962 1532
rect 1890 1513 1894 1515
rect 1890 1505 1894 1507
rect 1942 1514 1946 1516
rect 1942 1506 1946 1508
rect 1958 1513 1962 1515
rect 1958 1505 1962 1507
rect 1890 1488 1894 1490
rect 1890 1480 1894 1482
rect 1942 1489 1946 1491
rect 1942 1481 1946 1483
rect 1958 1488 1962 1490
rect 1958 1480 1962 1482
rect 1890 1463 1894 1465
rect 1890 1455 1894 1457
rect 1942 1464 1946 1466
rect 1942 1456 1946 1458
rect 1958 1463 1962 1465
rect 1958 1455 1962 1457
rect 1890 1438 1894 1440
rect 1890 1430 1894 1432
rect 1942 1439 1946 1441
rect 1942 1431 1946 1433
rect 1958 1438 1962 1440
rect 1958 1430 1962 1432
rect 1890 1413 1894 1415
rect 1890 1405 1894 1407
rect 1942 1414 1946 1416
rect 1942 1406 1946 1408
rect 1958 1413 1962 1415
rect 1958 1405 1962 1407
rect 1890 1388 1894 1390
rect 1890 1380 1894 1382
rect 1942 1389 1946 1391
rect 1942 1381 1946 1383
rect 1958 1388 1962 1390
rect 1758 1370 1760 1380
rect 1958 1380 1962 1382
rect 1890 1363 1894 1365
rect 1890 1355 1894 1357
rect 1942 1364 1946 1366
rect 1942 1356 1946 1358
rect 1958 1363 1962 1365
rect 1958 1355 1962 1357
rect 1890 1338 1894 1340
rect 1890 1330 1894 1332
rect 1942 1339 1946 1341
rect 1942 1331 1946 1333
rect 1958 1338 1962 1340
rect 1958 1330 1962 1332
rect 1890 1313 1894 1315
rect 1890 1305 1894 1307
rect 1942 1314 1946 1316
rect 1942 1306 1946 1308
rect 1958 1313 1962 1315
rect 1958 1305 1962 1307
rect 1890 1288 1894 1290
rect 1890 1280 1894 1282
rect 1942 1289 1946 1291
rect 1942 1281 1946 1283
rect 1958 1288 1962 1290
rect 1958 1280 1962 1282
rect 1890 1263 1894 1265
rect 1890 1255 1894 1257
rect 1942 1264 1946 1266
rect 1942 1256 1946 1258
rect 1958 1263 1962 1265
rect 1958 1255 1962 1257
rect 1890 1238 1894 1240
rect 1890 1230 1894 1232
rect 1942 1239 1946 1241
rect 1942 1231 1946 1233
rect 1958 1238 1962 1240
rect 1958 1230 1962 1232
rect 1890 1213 1894 1215
rect 1890 1205 1894 1207
rect 1942 1214 1946 1216
rect 1942 1206 1946 1208
rect 1958 1213 1962 1215
rect 912 1188 914 1198
rect 1958 1205 1962 1207
rect 1890 1188 1894 1190
rect 1890 1180 1894 1182
rect 1942 1189 1946 1191
rect 1942 1181 1946 1183
rect 1958 1188 1962 1190
rect 1958 1180 1962 1182
rect 1890 1163 1894 1165
rect 1890 1155 1894 1157
rect 1942 1164 1946 1166
rect 1942 1156 1946 1158
rect 1958 1163 1962 1165
rect 1958 1155 1962 1157
rect 1890 1138 1894 1140
rect 1890 1130 1894 1132
rect 1942 1139 1946 1141
rect 1942 1131 1946 1133
rect 1958 1138 1962 1140
rect 1958 1130 1962 1132
rect 1890 1113 1894 1115
rect 1890 1105 1894 1107
rect 1942 1114 1946 1116
rect 1942 1106 1946 1108
rect 1958 1113 1962 1115
rect 1958 1105 1962 1107
rect 1890 1088 1894 1090
rect 1890 1080 1894 1082
rect 1942 1089 1946 1091
rect 1942 1081 1946 1083
rect 1958 1088 1962 1090
rect 1958 1080 1962 1082
rect 1735 1055 1737 1065
rect 1753 1055 1755 1065
rect 1763 1055 1765 1065
rect 1890 1063 1894 1065
rect 1890 1055 1894 1057
rect 1942 1064 1946 1066
rect 1942 1056 1946 1058
rect 1958 1063 1962 1065
rect 1958 1055 1962 1057
rect 1890 1038 1894 1040
rect 1890 1030 1894 1032
rect 1942 1039 1946 1041
rect 1942 1031 1946 1033
rect 1958 1038 1962 1040
rect 1958 1030 1962 1032
rect 1890 1013 1894 1015
rect 1890 1005 1894 1007
rect 1942 1014 1946 1016
rect 1942 1006 1946 1008
rect 1958 1013 1962 1015
rect 1958 1005 1962 1007
rect 1890 988 1894 990
rect 1890 980 1894 982
rect 1942 989 1946 991
rect 1942 981 1946 983
rect 1958 988 1962 990
rect 1958 980 1962 982
rect 1890 963 1894 965
rect 1890 955 1894 957
rect 1942 964 1946 966
rect 1942 956 1946 958
rect 1958 963 1962 965
rect 1958 955 1962 957
rect 1890 938 1894 940
rect 1890 930 1894 932
rect 1942 939 1946 941
rect 1942 931 1946 933
rect 1958 938 1962 940
rect 1958 930 1962 932
rect 1890 913 1894 915
rect 1890 905 1894 907
rect 1942 914 1946 916
rect 1942 906 1946 908
rect 1958 913 1962 915
rect 1958 905 1962 907
rect 1890 888 1894 890
rect 1890 880 1894 882
rect 1942 889 1946 891
rect 1942 881 1946 883
rect 1958 888 1962 890
rect 1958 880 1962 882
rect 1890 863 1894 865
rect 1890 855 1894 857
rect 1942 864 1946 866
rect 1942 856 1946 858
rect 1958 863 1962 865
rect 1958 855 1962 857
rect 1890 838 1894 840
rect 1890 830 1894 832
rect 1942 839 1946 841
rect 1942 831 1946 833
rect 1958 838 1962 840
rect 1958 830 1962 832
rect 1890 813 1894 815
rect 1890 805 1894 807
rect 1942 814 1946 816
rect 1942 806 1946 808
rect 1958 813 1962 815
rect 1958 805 1962 807
rect 1890 788 1894 790
rect 1890 780 1894 782
rect 1942 789 1946 791
rect 1942 781 1946 783
rect 1958 788 1962 790
rect 1958 780 1962 782
rect 1890 763 1894 765
rect 1890 755 1894 757
rect 1942 764 1946 766
rect 1942 756 1946 758
rect 1958 763 1962 765
rect 1958 755 1962 757
rect 1890 738 1894 740
rect 1890 730 1894 732
rect 1942 739 1946 741
rect 1942 731 1946 733
rect 1958 738 1962 740
rect 1958 730 1962 732
rect 1890 713 1894 715
rect 1890 705 1894 707
rect 1942 714 1946 716
rect 1942 706 1946 708
rect 1958 713 1962 715
rect 1958 705 1962 707
rect 1890 688 1894 690
rect 1890 680 1894 682
rect 1942 689 1946 691
rect 1942 681 1946 683
rect 1958 688 1962 690
rect 1958 680 1962 682
rect 1890 663 1894 665
rect 1890 655 1894 657
rect 1942 664 1946 666
rect 1942 656 1946 658
rect 1958 663 1962 665
rect 1958 655 1962 657
rect 1890 638 1894 640
rect 1890 630 1894 632
rect 1942 639 1946 641
rect 1942 631 1946 633
rect 1958 638 1962 640
rect 1958 630 1962 632
rect 1890 613 1894 615
rect 1890 605 1894 607
rect 1942 614 1946 616
rect 1942 606 1946 608
rect 1958 613 1962 615
rect 1958 605 1962 607
rect 1890 588 1894 590
rect 1890 580 1894 582
rect 1942 589 1946 591
rect 1942 581 1946 583
rect 1958 588 1962 590
rect 1958 580 1962 582
rect 1890 563 1894 565
rect 1890 555 1894 557
rect 1942 564 1946 566
rect 1942 556 1946 558
rect 1958 563 1962 565
rect 1958 555 1962 557
rect 1890 538 1894 540
rect 1890 530 1894 532
rect 1942 539 1946 541
rect 1942 531 1946 533
rect 1958 538 1962 540
rect 1958 530 1962 532
rect 1890 513 1894 515
rect 1890 505 1894 507
rect 1942 514 1946 516
rect 1942 506 1946 508
rect 1958 513 1962 515
rect 1958 505 1962 507
rect 1890 488 1894 490
rect 1890 480 1894 482
rect 1942 489 1946 491
rect 1942 481 1946 483
rect 1958 488 1962 490
rect 1958 480 1962 482
rect 1890 463 1894 465
rect 1890 455 1894 457
rect 1942 464 1946 466
rect 1942 456 1946 458
rect 1958 463 1962 465
rect 1958 455 1962 457
rect 1890 438 1894 440
rect 1890 430 1894 432
rect 1942 439 1946 441
rect 1942 431 1946 433
rect 1958 438 1962 440
rect 1958 430 1962 432
rect 1890 413 1894 415
rect 1890 405 1894 407
rect 1942 414 1946 416
rect 1942 406 1946 408
rect 1958 413 1962 415
rect 1958 405 1962 407
rect 1890 388 1894 390
rect 1890 380 1894 382
rect 1942 389 1946 391
rect 1942 381 1946 383
rect 1958 388 1962 390
rect 1958 380 1962 382
rect 1890 363 1894 365
rect 1890 355 1894 357
rect 1942 364 1946 366
rect 1942 356 1946 358
rect 1958 363 1962 365
rect 1958 355 1962 357
rect 1890 338 1894 340
rect 1890 330 1894 332
rect 1942 339 1946 341
rect 1942 331 1946 333
rect 1958 338 1962 340
rect 1958 330 1962 332
rect 1890 313 1894 315
rect 1890 305 1894 307
rect 1942 314 1946 316
rect 1942 306 1946 308
rect 1958 313 1962 315
rect 1958 305 1962 307
rect 1890 288 1894 290
rect 1890 280 1894 282
rect 1942 289 1946 291
rect 1942 281 1946 283
rect 1958 288 1962 290
rect 1958 280 1962 282
rect 1890 263 1894 265
rect 1890 255 1894 257
rect 1942 264 1946 266
rect 1942 256 1946 258
rect 1958 263 1962 265
rect 1958 255 1962 257
rect 1890 238 1894 240
rect 1890 230 1894 232
rect 1942 239 1946 241
rect 1942 231 1946 233
rect 1958 238 1962 240
rect 1958 230 1962 232
rect 1890 213 1894 215
rect 1890 205 1894 207
rect 1942 214 1946 216
rect 1942 206 1946 208
rect 1958 213 1962 215
rect 1958 205 1962 207
rect 1890 188 1894 190
rect 1890 180 1894 182
rect 1942 189 1946 191
rect 1942 181 1946 183
rect 1958 188 1962 190
rect 1958 180 1962 182
rect 1890 163 1894 165
rect 1890 155 1894 157
rect 1942 164 1946 166
rect 1942 156 1946 158
rect 1958 163 1962 165
rect 1958 155 1962 157
rect 1890 138 1894 140
rect 1890 130 1894 132
rect 1942 139 1946 141
rect 1942 131 1946 133
rect 1958 138 1962 140
rect 1958 130 1962 132
rect 1890 113 1894 115
rect 1890 105 1894 107
rect 1942 114 1946 116
rect 1942 106 1946 108
rect 1958 113 1962 115
rect 1958 105 1962 107
rect 1890 88 1894 90
rect 1890 80 1894 82
rect 1942 89 1946 91
rect 1942 81 1946 83
rect 1958 88 1962 90
rect 1958 80 1962 82
rect 1890 63 1894 65
rect 1890 55 1894 57
rect 1942 64 1946 66
rect 1942 56 1946 58
rect 1958 63 1962 65
rect 1958 55 1962 57
rect 1890 38 1894 40
rect 1890 30 1894 32
rect 1942 39 1946 41
rect 1942 31 1946 33
rect 1958 38 1962 40
rect 1958 30 1962 32
<< ptransistor >>
rect 1904 2013 1912 2015
rect 1904 2005 1912 2007
rect 1924 2014 1932 2016
rect 1924 2006 1932 2008
rect 1972 2013 1980 2015
rect 1972 2005 1980 2007
rect 1904 1988 1912 1990
rect 1904 1980 1912 1982
rect 1924 1989 1932 1991
rect 1924 1981 1932 1983
rect 1972 1988 1980 1990
rect 1972 1980 1980 1982
rect 1904 1963 1912 1965
rect 1904 1955 1912 1957
rect 1924 1964 1932 1966
rect 1924 1956 1932 1958
rect 1972 1963 1980 1965
rect 1972 1955 1980 1957
rect 1904 1938 1912 1940
rect 1904 1930 1912 1932
rect 1924 1939 1932 1941
rect 1924 1931 1932 1933
rect 1972 1938 1980 1940
rect 1972 1930 1980 1932
rect 1904 1913 1912 1915
rect 1904 1905 1912 1907
rect 1924 1914 1932 1916
rect 1924 1906 1932 1908
rect 1972 1913 1980 1915
rect 1972 1905 1980 1907
rect 1904 1888 1912 1890
rect 1904 1880 1912 1882
rect 1924 1889 1932 1891
rect 1924 1881 1932 1883
rect 1972 1888 1980 1890
rect 1972 1880 1980 1882
rect 1904 1863 1912 1865
rect 1904 1855 1912 1857
rect 1924 1864 1932 1866
rect 1924 1856 1932 1858
rect 1972 1863 1980 1865
rect 1972 1855 1980 1857
rect 1904 1838 1912 1840
rect 1904 1830 1912 1832
rect 1924 1839 1932 1841
rect 1924 1831 1932 1833
rect 1972 1838 1980 1840
rect 1972 1830 1980 1832
rect 1904 1813 1912 1815
rect 1904 1805 1912 1807
rect 1924 1814 1932 1816
rect 1924 1806 1932 1808
rect 1972 1813 1980 1815
rect 1972 1805 1980 1807
rect 1904 1788 1912 1790
rect 1904 1780 1912 1782
rect 1924 1789 1932 1791
rect 1924 1781 1932 1783
rect 1972 1788 1980 1790
rect 1972 1780 1980 1782
rect 1904 1763 1912 1765
rect 1904 1755 1912 1757
rect 1924 1764 1932 1766
rect 1924 1756 1932 1758
rect 1972 1763 1980 1765
rect 1972 1755 1980 1757
rect 1904 1738 1912 1740
rect 1904 1730 1912 1732
rect 1924 1739 1932 1741
rect 1924 1731 1932 1733
rect 1972 1738 1980 1740
rect 1972 1730 1980 1732
rect 1904 1713 1912 1715
rect 1904 1705 1912 1707
rect 1924 1714 1932 1716
rect 1924 1706 1932 1708
rect 1972 1713 1980 1715
rect 1972 1705 1980 1707
rect 1904 1688 1912 1690
rect 1904 1680 1912 1682
rect 1924 1689 1932 1691
rect 1924 1681 1932 1683
rect 1972 1688 1980 1690
rect 1972 1680 1980 1682
rect 1904 1663 1912 1665
rect 1904 1655 1912 1657
rect 1924 1664 1932 1666
rect 1924 1656 1932 1658
rect 1972 1663 1980 1665
rect 1972 1655 1980 1657
rect 1904 1638 1912 1640
rect 1904 1630 1912 1632
rect 1924 1639 1932 1641
rect 1924 1631 1932 1633
rect 1972 1638 1980 1640
rect 1972 1630 1980 1632
rect 1904 1613 1912 1615
rect 1904 1605 1912 1607
rect 1924 1614 1932 1616
rect 1924 1606 1932 1608
rect 1972 1613 1980 1615
rect 1972 1605 1980 1607
rect 1904 1588 1912 1590
rect 1904 1580 1912 1582
rect 1924 1589 1932 1591
rect 1924 1581 1932 1583
rect 1972 1588 1980 1590
rect 1972 1580 1980 1582
rect 1904 1563 1912 1565
rect 1904 1555 1912 1557
rect 1924 1564 1932 1566
rect 1924 1556 1932 1558
rect 1972 1563 1980 1565
rect 1972 1555 1980 1557
rect 1904 1538 1912 1540
rect 1904 1530 1912 1532
rect 1924 1539 1932 1541
rect 1924 1531 1932 1533
rect 1972 1538 1980 1540
rect 1972 1530 1980 1532
rect 1904 1513 1912 1515
rect 1904 1505 1912 1507
rect 1924 1514 1932 1516
rect 1924 1506 1932 1508
rect 1972 1513 1980 1515
rect 1972 1505 1980 1507
rect 1904 1488 1912 1490
rect 1904 1480 1912 1482
rect 1924 1489 1932 1491
rect 1924 1481 1932 1483
rect 1972 1488 1980 1490
rect 1972 1480 1980 1482
rect 1904 1463 1912 1465
rect 1904 1455 1912 1457
rect 1924 1464 1932 1466
rect 1924 1456 1932 1458
rect 1972 1463 1980 1465
rect 1972 1455 1980 1457
rect 1904 1438 1912 1440
rect 1904 1430 1912 1432
rect 1924 1439 1932 1441
rect 1924 1431 1932 1433
rect 1972 1438 1980 1440
rect 1972 1430 1980 1432
rect 1758 1390 1760 1410
rect 1904 1413 1912 1415
rect 1904 1405 1912 1407
rect 1924 1414 1932 1416
rect 1924 1406 1932 1408
rect 1972 1413 1980 1415
rect 1972 1405 1980 1407
rect 1904 1388 1912 1390
rect 1904 1380 1912 1382
rect 1924 1389 1932 1391
rect 1924 1381 1932 1383
rect 1972 1388 1980 1390
rect 1972 1380 1980 1382
rect 1904 1363 1912 1365
rect 1904 1355 1912 1357
rect 1924 1364 1932 1366
rect 1924 1356 1932 1358
rect 1972 1363 1980 1365
rect 1972 1355 1980 1357
rect 1904 1338 1912 1340
rect 1904 1330 1912 1332
rect 1924 1339 1932 1341
rect 1924 1331 1932 1333
rect 1972 1338 1980 1340
rect 1972 1330 1980 1332
rect 1904 1313 1912 1315
rect 1904 1305 1912 1307
rect 1924 1314 1932 1316
rect 1924 1306 1932 1308
rect 1972 1313 1980 1315
rect 1972 1305 1980 1307
rect 1904 1288 1912 1290
rect 1904 1280 1912 1282
rect 1924 1289 1932 1291
rect 1924 1281 1932 1283
rect 1972 1288 1980 1290
rect 1972 1280 1980 1282
rect 1904 1263 1912 1265
rect 1904 1255 1912 1257
rect 1924 1264 1932 1266
rect 1924 1256 1932 1258
rect 1972 1263 1980 1265
rect 1972 1255 1980 1257
rect 1904 1238 1912 1240
rect 1904 1230 1912 1232
rect 1924 1239 1932 1241
rect 1924 1231 1932 1233
rect 1972 1238 1980 1240
rect 1972 1230 1980 1232
rect 1904 1213 1912 1215
rect 1904 1205 1912 1207
rect 1924 1214 1932 1216
rect 1924 1206 1932 1208
rect 1972 1213 1980 1215
rect 1972 1205 1980 1207
rect 1904 1188 1912 1190
rect 1904 1180 1912 1182
rect 1924 1189 1932 1191
rect 1924 1181 1932 1183
rect 1972 1188 1980 1190
rect 912 1158 914 1178
rect 1972 1180 1980 1182
rect 1904 1163 1912 1165
rect 1904 1155 1912 1157
rect 1924 1164 1932 1166
rect 1924 1156 1932 1158
rect 1972 1163 1980 1165
rect 1972 1155 1980 1157
rect 1904 1138 1912 1140
rect 1904 1130 1912 1132
rect 1924 1139 1932 1141
rect 1924 1131 1932 1133
rect 1972 1138 1980 1140
rect 1972 1130 1980 1132
rect 1904 1113 1912 1115
rect 1904 1105 1912 1107
rect 1924 1114 1932 1116
rect 1924 1106 1932 1108
rect 1972 1113 1980 1115
rect 1735 1075 1737 1093
rect 1753 1075 1755 1093
rect 1763 1075 1765 1093
rect 1972 1105 1980 1107
rect 1904 1088 1912 1090
rect 1904 1080 1912 1082
rect 1924 1089 1932 1091
rect 1924 1081 1932 1083
rect 1972 1088 1980 1090
rect 1972 1080 1980 1082
rect 1904 1063 1912 1065
rect 1904 1055 1912 1057
rect 1924 1064 1932 1066
rect 1924 1056 1932 1058
rect 1972 1063 1980 1065
rect 1972 1055 1980 1057
rect 1904 1038 1912 1040
rect 1904 1030 1912 1032
rect 1924 1039 1932 1041
rect 1924 1031 1932 1033
rect 1972 1038 1980 1040
rect 1972 1030 1980 1032
rect 1904 1013 1912 1015
rect 1904 1005 1912 1007
rect 1924 1014 1932 1016
rect 1924 1006 1932 1008
rect 1972 1013 1980 1015
rect 1972 1005 1980 1007
rect 1904 988 1912 990
rect 1904 980 1912 982
rect 1924 989 1932 991
rect 1924 981 1932 983
rect 1972 988 1980 990
rect 1972 980 1980 982
rect 1904 963 1912 965
rect 1904 955 1912 957
rect 1924 964 1932 966
rect 1924 956 1932 958
rect 1972 963 1980 965
rect 1972 955 1980 957
rect 1904 938 1912 940
rect 1904 930 1912 932
rect 1924 939 1932 941
rect 1924 931 1932 933
rect 1972 938 1980 940
rect 1972 930 1980 932
rect 1904 913 1912 915
rect 1904 905 1912 907
rect 1924 914 1932 916
rect 1924 906 1932 908
rect 1972 913 1980 915
rect 1972 905 1980 907
rect 1904 888 1912 890
rect 1904 880 1912 882
rect 1924 889 1932 891
rect 1924 881 1932 883
rect 1972 888 1980 890
rect 1972 880 1980 882
rect 1904 863 1912 865
rect 1904 855 1912 857
rect 1924 864 1932 866
rect 1924 856 1932 858
rect 1972 863 1980 865
rect 1972 855 1980 857
rect 1904 838 1912 840
rect 1904 830 1912 832
rect 1924 839 1932 841
rect 1924 831 1932 833
rect 1972 838 1980 840
rect 1972 830 1980 832
rect 1904 813 1912 815
rect 1904 805 1912 807
rect 1924 814 1932 816
rect 1924 806 1932 808
rect 1972 813 1980 815
rect 1972 805 1980 807
rect 1904 788 1912 790
rect 1904 780 1912 782
rect 1924 789 1932 791
rect 1924 781 1932 783
rect 1972 788 1980 790
rect 1972 780 1980 782
rect 1904 763 1912 765
rect 1904 755 1912 757
rect 1924 764 1932 766
rect 1924 756 1932 758
rect 1972 763 1980 765
rect 1972 755 1980 757
rect 1904 738 1912 740
rect 1904 730 1912 732
rect 1924 739 1932 741
rect 1924 731 1932 733
rect 1972 738 1980 740
rect 1972 730 1980 732
rect 1904 713 1912 715
rect 1904 705 1912 707
rect 1924 714 1932 716
rect 1924 706 1932 708
rect 1972 713 1980 715
rect 1972 705 1980 707
rect 1904 688 1912 690
rect 1904 680 1912 682
rect 1924 689 1932 691
rect 1924 681 1932 683
rect 1972 688 1980 690
rect 1972 680 1980 682
rect 1904 663 1912 665
rect 1904 655 1912 657
rect 1924 664 1932 666
rect 1924 656 1932 658
rect 1972 663 1980 665
rect 1972 655 1980 657
rect 1904 638 1912 640
rect 1904 630 1912 632
rect 1924 639 1932 641
rect 1924 631 1932 633
rect 1972 638 1980 640
rect 1972 630 1980 632
rect 1904 613 1912 615
rect 1904 605 1912 607
rect 1924 614 1932 616
rect 1924 606 1932 608
rect 1972 613 1980 615
rect 1972 605 1980 607
rect 1904 588 1912 590
rect 1904 580 1912 582
rect 1924 589 1932 591
rect 1924 581 1932 583
rect 1972 588 1980 590
rect 1972 580 1980 582
rect 1904 563 1912 565
rect 1904 555 1912 557
rect 1924 564 1932 566
rect 1924 556 1932 558
rect 1972 563 1980 565
rect 1972 555 1980 557
rect 1904 538 1912 540
rect 1904 530 1912 532
rect 1924 539 1932 541
rect 1924 531 1932 533
rect 1972 538 1980 540
rect 1972 530 1980 532
rect 1904 513 1912 515
rect 1904 505 1912 507
rect 1924 514 1932 516
rect 1924 506 1932 508
rect 1972 513 1980 515
rect 1972 505 1980 507
rect 1904 488 1912 490
rect 1904 480 1912 482
rect 1924 489 1932 491
rect 1924 481 1932 483
rect 1972 488 1980 490
rect 1972 480 1980 482
rect 1904 463 1912 465
rect 1904 455 1912 457
rect 1924 464 1932 466
rect 1924 456 1932 458
rect 1972 463 1980 465
rect 1972 455 1980 457
rect 1904 438 1912 440
rect 1904 430 1912 432
rect 1924 439 1932 441
rect 1924 431 1932 433
rect 1972 438 1980 440
rect 1972 430 1980 432
rect 1904 413 1912 415
rect 1904 405 1912 407
rect 1924 414 1932 416
rect 1924 406 1932 408
rect 1972 413 1980 415
rect 1972 405 1980 407
rect 1904 388 1912 390
rect 1904 380 1912 382
rect 1924 389 1932 391
rect 1924 381 1932 383
rect 1972 388 1980 390
rect 1972 380 1980 382
rect 1904 363 1912 365
rect 1904 355 1912 357
rect 1924 364 1932 366
rect 1924 356 1932 358
rect 1972 363 1980 365
rect 1972 355 1980 357
rect 1904 338 1912 340
rect 1904 330 1912 332
rect 1924 339 1932 341
rect 1924 331 1932 333
rect 1972 338 1980 340
rect 1972 330 1980 332
rect 1904 313 1912 315
rect 1904 305 1912 307
rect 1924 314 1932 316
rect 1924 306 1932 308
rect 1972 313 1980 315
rect 1972 305 1980 307
rect 1904 288 1912 290
rect 1904 280 1912 282
rect 1924 289 1932 291
rect 1924 281 1932 283
rect 1972 288 1980 290
rect 1972 280 1980 282
rect 1904 263 1912 265
rect 1904 255 1912 257
rect 1924 264 1932 266
rect 1924 256 1932 258
rect 1972 263 1980 265
rect 1972 255 1980 257
rect 1904 238 1912 240
rect 1904 230 1912 232
rect 1924 239 1932 241
rect 1924 231 1932 233
rect 1972 238 1980 240
rect 1972 230 1980 232
rect 1904 213 1912 215
rect 1904 205 1912 207
rect 1924 214 1932 216
rect 1924 206 1932 208
rect 1972 213 1980 215
rect 1972 205 1980 207
rect 1904 188 1912 190
rect 1904 180 1912 182
rect 1924 189 1932 191
rect 1924 181 1932 183
rect 1972 188 1980 190
rect 1972 180 1980 182
rect 1904 163 1912 165
rect 1904 155 1912 157
rect 1924 164 1932 166
rect 1924 156 1932 158
rect 1972 163 1980 165
rect 1972 155 1980 157
rect 1904 138 1912 140
rect 1904 130 1912 132
rect 1924 139 1932 141
rect 1924 131 1932 133
rect 1972 138 1980 140
rect 1972 130 1980 132
rect 1904 113 1912 115
rect 1904 105 1912 107
rect 1924 114 1932 116
rect 1924 106 1932 108
rect 1972 113 1980 115
rect 1972 105 1980 107
rect 1904 88 1912 90
rect 1904 80 1912 82
rect 1924 89 1932 91
rect 1924 81 1932 83
rect 1972 88 1980 90
rect 1972 80 1980 82
rect 1904 63 1912 65
rect 1904 55 1912 57
rect 1924 64 1932 66
rect 1924 56 1932 58
rect 1972 63 1980 65
rect 1972 55 1980 57
rect 1904 38 1912 40
rect 1904 30 1912 32
rect 1924 39 1932 41
rect 1924 31 1932 33
rect 1972 38 1980 40
rect 1972 30 1980 32
<< polycontact >>
rect 1867 2019 1874 2026
rect 1935 2019 1939 2023
rect 1897 2006 1901 2010
rect 1935 2011 1939 2015
rect 1897 1998 1901 2002
rect 1965 2006 1969 2010
rect 1935 1994 1939 1998
rect 1965 1998 1969 2002
rect 1897 1981 1901 1985
rect 1935 1986 1939 1990
rect 1897 1973 1901 1977
rect 1965 1981 1969 1985
rect 1935 1969 1939 1973
rect 1965 1973 1969 1977
rect 1897 1956 1901 1960
rect 1935 1961 1939 1965
rect 1897 1948 1901 1952
rect 1965 1956 1969 1960
rect 1935 1944 1939 1948
rect 1965 1948 1969 1952
rect 1897 1931 1901 1935
rect 1935 1936 1939 1940
rect 1897 1923 1901 1927
rect 1965 1931 1969 1935
rect 1935 1919 1939 1923
rect 1965 1923 1969 1927
rect 1897 1906 1901 1910
rect 1935 1911 1939 1915
rect 1897 1898 1901 1902
rect 1965 1906 1969 1910
rect 1935 1894 1939 1898
rect 1965 1898 1969 1902
rect 1897 1881 1901 1885
rect 1935 1886 1939 1890
rect 1897 1873 1901 1877
rect 1965 1881 1969 1885
rect 1935 1869 1939 1873
rect 1965 1873 1969 1877
rect 1897 1856 1901 1860
rect 1935 1861 1939 1865
rect 1897 1848 1901 1852
rect 1965 1856 1969 1860
rect 1935 1844 1939 1848
rect 1965 1848 1969 1852
rect 1897 1831 1901 1835
rect 1935 1836 1939 1840
rect 1897 1823 1901 1827
rect 1965 1831 1969 1835
rect 1935 1819 1939 1823
rect 1965 1823 1969 1827
rect 1897 1806 1901 1810
rect 1935 1811 1939 1815
rect 1897 1798 1901 1802
rect 1965 1806 1969 1810
rect 1935 1794 1939 1798
rect 1965 1798 1969 1802
rect 1897 1781 1901 1785
rect 1935 1786 1939 1790
rect 1897 1773 1901 1777
rect 1965 1781 1969 1785
rect 1935 1769 1939 1773
rect 1965 1773 1969 1777
rect 1897 1756 1901 1760
rect 1935 1761 1939 1765
rect 1897 1748 1901 1752
rect 1965 1756 1969 1760
rect 1935 1744 1939 1748
rect 1965 1748 1969 1752
rect 1897 1731 1901 1735
rect 1935 1736 1939 1740
rect 1897 1723 1901 1727
rect 1965 1731 1969 1735
rect 1935 1719 1939 1723
rect 1965 1723 1969 1727
rect 1897 1706 1901 1710
rect 1935 1711 1939 1715
rect 1897 1698 1901 1702
rect 1965 1706 1969 1710
rect 1935 1694 1939 1698
rect 1965 1698 1969 1702
rect 1897 1681 1901 1685
rect 1935 1686 1939 1690
rect 1897 1673 1901 1677
rect 1424 1664 1430 1670
rect 1965 1681 1969 1685
rect 1935 1669 1939 1673
rect 1965 1673 1969 1677
rect 1897 1656 1901 1660
rect 1935 1661 1939 1665
rect 1897 1648 1901 1652
rect 910 1635 915 1643
rect 1965 1656 1969 1660
rect 1935 1644 1939 1648
rect 1965 1648 1969 1652
rect 1897 1631 1901 1635
rect 1935 1636 1939 1640
rect 1897 1623 1901 1627
rect 1965 1631 1969 1635
rect 1935 1619 1939 1623
rect 1965 1623 1969 1627
rect 1897 1606 1901 1610
rect 1935 1611 1939 1615
rect 1897 1598 1901 1602
rect 1965 1606 1969 1610
rect 1935 1594 1939 1598
rect 1965 1598 1969 1602
rect 1897 1581 1901 1585
rect 1935 1586 1939 1590
rect 1897 1573 1901 1577
rect 1965 1581 1969 1585
rect 1935 1569 1939 1573
rect 1965 1573 1969 1577
rect 1897 1556 1901 1560
rect 1935 1561 1939 1565
rect 1897 1548 1901 1552
rect 1965 1556 1969 1560
rect 1935 1544 1939 1548
rect 1965 1548 1969 1552
rect 1897 1531 1901 1535
rect 1935 1536 1939 1540
rect 1897 1523 1901 1527
rect 1965 1531 1969 1535
rect 1935 1519 1939 1523
rect 1965 1523 1969 1527
rect 1897 1506 1901 1510
rect 1935 1511 1939 1515
rect 1897 1498 1901 1502
rect 1965 1506 1969 1510
rect 1935 1494 1939 1498
rect 1965 1498 1969 1502
rect 1897 1481 1901 1485
rect 1935 1486 1939 1490
rect 1897 1473 1901 1477
rect 1965 1481 1969 1485
rect 1935 1469 1939 1473
rect 1965 1473 1969 1477
rect 1897 1456 1901 1460
rect 1935 1461 1939 1465
rect 1897 1448 1901 1452
rect 1707 1434 1715 1442
rect 1965 1456 1969 1460
rect 1935 1444 1939 1448
rect 1965 1448 1969 1452
rect 1897 1431 1901 1435
rect 1935 1436 1939 1440
rect 1897 1423 1901 1427
rect 1965 1431 1969 1435
rect 1935 1419 1939 1423
rect 1965 1423 1969 1427
rect 1897 1406 1901 1410
rect 1935 1411 1939 1415
rect 1897 1398 1901 1402
rect 1965 1406 1969 1410
rect 1935 1394 1939 1398
rect 1965 1398 1969 1402
rect 1787 1383 1792 1387
rect 1897 1381 1901 1385
rect 1935 1386 1939 1390
rect 1897 1373 1901 1377
rect 1965 1381 1969 1385
rect 1935 1369 1939 1373
rect 1965 1373 1969 1377
rect 1897 1356 1901 1360
rect 1935 1361 1939 1365
rect 1897 1348 1901 1352
rect 1965 1356 1969 1360
rect 1935 1344 1939 1348
rect 1965 1348 1969 1352
rect 1897 1331 1901 1335
rect 1935 1336 1939 1340
rect 1897 1323 1901 1327
rect 1965 1331 1969 1335
rect 1935 1319 1939 1323
rect 1965 1323 1969 1327
rect 1897 1306 1901 1310
rect 1935 1311 1939 1315
rect 1897 1298 1901 1302
rect 1965 1306 1969 1310
rect 1935 1294 1939 1298
rect 1965 1298 1969 1302
rect 1897 1281 1901 1285
rect 1935 1286 1939 1290
rect 1897 1273 1901 1277
rect 1965 1281 1969 1285
rect 1935 1269 1939 1273
rect 1965 1273 1969 1277
rect 1897 1256 1901 1260
rect 1935 1261 1939 1265
rect 1897 1248 1901 1252
rect 1965 1256 1969 1260
rect 1935 1244 1939 1248
rect 1965 1248 1969 1252
rect 1897 1231 1901 1235
rect 1935 1236 1939 1240
rect 1897 1223 1901 1227
rect 1965 1231 1969 1235
rect 1935 1219 1939 1223
rect 1965 1223 1969 1227
rect 1897 1206 1901 1210
rect 1935 1211 1939 1215
rect 1897 1198 1901 1202
rect 1965 1206 1969 1210
rect 1935 1194 1939 1198
rect 1965 1198 1969 1202
rect 914 1181 918 1185
rect 1897 1181 1901 1185
rect 1935 1186 1939 1190
rect 1897 1173 1901 1177
rect 1965 1181 1969 1185
rect 1935 1169 1939 1173
rect 1965 1173 1969 1177
rect 1897 1156 1901 1160
rect 1935 1161 1939 1165
rect 1897 1148 1901 1152
rect 1965 1156 1969 1160
rect 1935 1144 1939 1148
rect 1965 1148 1969 1152
rect 1897 1131 1901 1135
rect 1935 1136 1939 1140
rect 1897 1123 1901 1127
rect 1965 1131 1969 1135
rect 1935 1119 1939 1123
rect 1965 1123 1969 1127
rect 1897 1106 1901 1110
rect 1935 1111 1939 1115
rect 1750 1097 1754 1101
rect 1764 1097 1768 1101
rect 1897 1098 1901 1102
rect 1965 1106 1969 1110
rect 1935 1094 1939 1098
rect 1965 1098 1969 1102
rect 1897 1081 1901 1085
rect 1935 1086 1939 1090
rect 1736 1068 1740 1072
rect 1897 1073 1901 1077
rect 1965 1081 1969 1085
rect 1935 1069 1939 1073
rect 1965 1073 1969 1077
rect 1897 1056 1901 1060
rect 1935 1061 1939 1065
rect 1897 1048 1901 1052
rect 1965 1056 1969 1060
rect 1935 1044 1939 1048
rect 1965 1048 1969 1052
rect 1897 1031 1901 1035
rect 1935 1036 1939 1040
rect 1897 1023 1901 1027
rect 1965 1031 1969 1035
rect 1935 1019 1939 1023
rect 1965 1023 1969 1027
rect 1897 1006 1901 1010
rect 1935 1011 1939 1015
rect 1897 998 1901 1002
rect 1965 1006 1969 1010
rect 1935 994 1939 998
rect 1965 998 1969 1002
rect 1897 981 1901 985
rect 1935 986 1939 990
rect 1897 973 1901 977
rect 1965 981 1969 985
rect 1935 969 1939 973
rect 1965 973 1969 977
rect 1897 956 1901 960
rect 1935 961 1939 965
rect 1897 948 1901 952
rect 1965 956 1969 960
rect 1935 944 1939 948
rect 1965 948 1969 952
rect 1897 931 1901 935
rect 1935 936 1939 940
rect 1897 923 1901 927
rect 1965 931 1969 935
rect 1935 919 1939 923
rect 1965 923 1969 927
rect 1897 906 1901 910
rect 1935 911 1939 915
rect 1897 898 1901 902
rect 1965 906 1969 910
rect 1935 894 1939 898
rect 1965 898 1969 902
rect 1897 881 1901 885
rect 1935 886 1939 890
rect 1897 873 1901 877
rect 1965 881 1969 885
rect 1935 869 1939 873
rect 1965 873 1969 877
rect 1897 856 1901 860
rect 1935 861 1939 865
rect 1897 848 1901 852
rect 1965 856 1969 860
rect 1935 844 1939 848
rect 1965 848 1969 852
rect 1897 831 1901 835
rect 1935 836 1939 840
rect 1897 823 1901 827
rect 1965 831 1969 835
rect 1935 819 1939 823
rect 1965 823 1969 827
rect 1897 806 1901 810
rect 1935 811 1939 815
rect 1897 798 1901 802
rect 1965 806 1969 810
rect 1935 794 1939 798
rect 1965 798 1969 802
rect 1897 781 1901 785
rect 1935 786 1939 790
rect 1897 773 1901 777
rect 1965 781 1969 785
rect 1935 769 1939 773
rect 1965 773 1969 777
rect 1897 756 1901 760
rect 1935 761 1939 765
rect 1790 745 1795 753
rect 1897 748 1901 752
rect 1965 756 1969 760
rect 1935 744 1939 748
rect 1965 748 1969 752
rect 1897 731 1901 735
rect 1935 736 1939 740
rect 1897 723 1901 727
rect 1965 731 1969 735
rect 1935 719 1939 723
rect 1965 723 1969 727
rect 1897 706 1901 710
rect 1935 711 1939 715
rect 1897 698 1901 702
rect 1965 706 1969 710
rect 1935 694 1939 698
rect 1965 698 1969 702
rect 1897 681 1901 685
rect 1935 686 1939 690
rect 1897 673 1901 677
rect 1965 681 1969 685
rect 1935 669 1939 673
rect 1965 673 1969 677
rect 1897 656 1901 660
rect 1935 661 1939 665
rect 1897 648 1901 652
rect 1965 656 1969 660
rect 1935 644 1939 648
rect 1965 648 1969 652
rect 1897 631 1901 635
rect 1935 636 1939 640
rect 1897 623 1901 627
rect 1965 631 1969 635
rect 1935 619 1939 623
rect 1965 623 1969 627
rect 1897 606 1901 610
rect 1935 611 1939 615
rect 1897 598 1901 602
rect 1965 606 1969 610
rect 1935 594 1939 598
rect 1965 598 1969 602
rect 1897 581 1901 585
rect 1935 586 1939 590
rect 1897 573 1901 577
rect 1965 581 1969 585
rect 1935 569 1939 573
rect 1965 573 1969 577
rect 1897 556 1901 560
rect 1935 561 1939 565
rect 1897 548 1901 552
rect 1965 556 1969 560
rect 1935 544 1939 548
rect 1965 548 1969 552
rect 1897 531 1901 535
rect 1935 536 1939 540
rect 1897 523 1901 527
rect 1965 531 1969 535
rect 1935 519 1939 523
rect 1965 523 1969 527
rect 1897 506 1901 510
rect 1935 511 1939 515
rect 1897 498 1901 502
rect 1965 506 1969 510
rect 1935 494 1939 498
rect 1965 498 1969 502
rect 1897 481 1901 485
rect 1935 486 1939 490
rect 1897 473 1901 477
rect 1965 481 1969 485
rect 1935 469 1939 473
rect 1965 473 1969 477
rect 1897 456 1901 460
rect 1935 461 1939 465
rect 1897 448 1901 452
rect 1965 456 1969 460
rect 1935 444 1939 448
rect 1965 448 1969 452
rect 1897 431 1901 435
rect 1935 436 1939 440
rect 1897 423 1901 427
rect 1965 431 1969 435
rect 1935 419 1939 423
rect 1965 423 1969 427
rect 1897 406 1901 410
rect 1935 411 1939 415
rect 1897 398 1901 402
rect 1965 406 1969 410
rect 1935 394 1939 398
rect 1965 398 1969 402
rect 1897 381 1901 385
rect 1935 386 1939 390
rect 1897 373 1901 377
rect 1965 381 1969 385
rect 1935 369 1939 373
rect 1965 373 1969 377
rect 1897 356 1901 360
rect 1935 361 1939 365
rect 1897 348 1901 352
rect 1965 356 1969 360
rect 1935 344 1939 348
rect 1965 348 1969 352
rect 1897 331 1901 335
rect 1935 336 1939 340
rect 1897 323 1901 327
rect 1965 331 1969 335
rect 1935 319 1939 323
rect 1965 323 1969 327
rect 1897 306 1901 310
rect 1935 311 1939 315
rect 1897 298 1901 302
rect 1965 306 1969 310
rect 1935 294 1939 298
rect 1965 298 1969 302
rect 1897 281 1901 285
rect 1935 286 1939 290
rect 1897 273 1901 277
rect 1965 281 1969 285
rect 1935 269 1939 273
rect 1965 273 1969 277
rect 1897 256 1901 260
rect 1935 261 1939 265
rect 1897 248 1901 252
rect 1965 256 1969 260
rect 1935 244 1939 248
rect 1965 248 1969 252
rect 1897 231 1901 235
rect 1935 236 1939 240
rect 1897 223 1901 227
rect 1965 231 1969 235
rect 1935 219 1939 223
rect 1965 223 1969 227
rect 1897 206 1901 210
rect 1935 211 1939 215
rect 1897 198 1901 202
rect 1965 206 1969 210
rect 1935 194 1939 198
rect 1965 198 1969 202
rect 1897 181 1901 185
rect 1935 186 1939 190
rect 1897 173 1901 177
rect 1965 181 1969 185
rect 1935 169 1939 173
rect 1965 173 1969 177
rect 1897 156 1901 160
rect 1935 161 1939 165
rect 1897 148 1901 152
rect 1965 156 1969 160
rect 1935 144 1939 148
rect 1965 148 1969 152
rect 1897 131 1901 135
rect 1935 136 1939 140
rect 1897 123 1901 127
rect 1965 131 1969 135
rect 1935 119 1939 123
rect 1965 123 1969 127
rect 1897 106 1901 110
rect 1935 111 1939 115
rect 1897 98 1901 102
rect 1965 106 1969 110
rect 1935 94 1939 98
rect 1965 98 1969 102
rect 1897 81 1901 85
rect 1935 86 1939 90
rect 1897 73 1901 77
rect 1965 81 1969 85
rect 1935 69 1939 73
rect 1965 73 1969 77
rect 1897 56 1901 60
rect 1935 61 1939 65
rect 1897 48 1901 52
rect 1965 56 1969 60
rect 1935 44 1939 48
rect 1965 48 1969 52
rect 1897 31 1901 35
rect 1935 36 1939 40
rect 1897 23 1901 27
rect 1965 31 1969 35
rect 1965 23 1969 27
rect 1801 17 1807 23
<< ndcontact >>
rect 1890 2016 1894 2020
rect 1942 2017 1946 2021
rect 1958 2016 1962 2020
rect 1890 2008 1894 2012
rect 1942 2009 1946 2013
rect 1958 2008 1962 2012
rect 1890 2000 1894 2004
rect 1890 1991 1894 1995
rect 1942 2001 1946 2005
rect 1958 2000 1962 2004
rect 1942 1992 1946 1996
rect 1958 1991 1962 1995
rect 1890 1983 1894 1987
rect 1942 1984 1946 1988
rect 1958 1983 1962 1987
rect 1890 1975 1894 1979
rect 1890 1966 1894 1970
rect 1942 1976 1946 1980
rect 1958 1975 1962 1979
rect 1942 1967 1946 1971
rect 1958 1966 1962 1970
rect 1890 1958 1894 1962
rect 1942 1959 1946 1963
rect 1958 1958 1962 1962
rect 1890 1950 1894 1954
rect 1890 1941 1894 1945
rect 1942 1951 1946 1955
rect 1958 1950 1962 1954
rect 1942 1942 1946 1946
rect 1958 1941 1962 1945
rect 1890 1933 1894 1937
rect 1942 1934 1946 1938
rect 1958 1933 1962 1937
rect 1890 1925 1894 1929
rect 1890 1916 1894 1920
rect 1942 1926 1946 1930
rect 1958 1925 1962 1929
rect 1942 1917 1946 1921
rect 1958 1916 1962 1920
rect 1890 1908 1894 1912
rect 1942 1909 1946 1913
rect 1958 1908 1962 1912
rect 1890 1900 1894 1904
rect 1890 1891 1894 1895
rect 1942 1901 1946 1905
rect 1958 1900 1962 1904
rect 1942 1892 1946 1896
rect 1958 1891 1962 1895
rect 1890 1883 1894 1887
rect 1942 1884 1946 1888
rect 1958 1883 1962 1887
rect 1890 1875 1894 1879
rect 1890 1866 1894 1870
rect 1942 1876 1946 1880
rect 1958 1875 1962 1879
rect 1942 1867 1946 1871
rect 1958 1866 1962 1870
rect 1890 1858 1894 1862
rect 1942 1859 1946 1863
rect 1958 1858 1962 1862
rect 1890 1850 1894 1854
rect 1890 1841 1894 1845
rect 1942 1851 1946 1855
rect 1958 1850 1962 1854
rect 1942 1842 1946 1846
rect 1958 1841 1962 1845
rect 1890 1833 1894 1837
rect 1942 1834 1946 1838
rect 1958 1833 1962 1837
rect 1890 1825 1894 1829
rect 1890 1816 1894 1820
rect 1942 1826 1946 1830
rect 1958 1825 1962 1829
rect 1942 1817 1946 1821
rect 1958 1816 1962 1820
rect 1890 1808 1894 1812
rect 1942 1809 1946 1813
rect 1958 1808 1962 1812
rect 1890 1800 1894 1804
rect 1890 1791 1894 1795
rect 1942 1801 1946 1805
rect 1958 1800 1962 1804
rect 1942 1792 1946 1796
rect 1958 1791 1962 1795
rect 1890 1783 1894 1787
rect 1942 1784 1946 1788
rect 1958 1783 1962 1787
rect 1890 1775 1894 1779
rect 1890 1766 1894 1770
rect 1942 1776 1946 1780
rect 1958 1775 1962 1779
rect 1942 1767 1946 1771
rect 1958 1766 1962 1770
rect 1890 1758 1894 1762
rect 1942 1759 1946 1763
rect 1958 1758 1962 1762
rect 1890 1750 1894 1754
rect 1890 1741 1894 1745
rect 1942 1751 1946 1755
rect 1958 1750 1962 1754
rect 1942 1742 1946 1746
rect 1958 1741 1962 1745
rect 1890 1733 1894 1737
rect 1942 1734 1946 1738
rect 1958 1733 1962 1737
rect 1890 1725 1894 1729
rect 1890 1716 1894 1720
rect 1942 1726 1946 1730
rect 1958 1725 1962 1729
rect 1942 1717 1946 1721
rect 1958 1716 1962 1720
rect 1890 1708 1894 1712
rect 1942 1709 1946 1713
rect 1958 1708 1962 1712
rect 1890 1700 1894 1704
rect 1890 1691 1894 1695
rect 1942 1701 1946 1705
rect 1958 1700 1962 1704
rect 1942 1692 1946 1696
rect 1958 1691 1962 1695
rect 1890 1683 1894 1687
rect 1942 1684 1946 1688
rect 1958 1683 1962 1687
rect 1890 1675 1894 1679
rect 1890 1666 1894 1670
rect 1942 1676 1946 1680
rect 1958 1675 1962 1679
rect 1942 1667 1946 1671
rect 1958 1666 1962 1670
rect 1890 1658 1894 1662
rect 1942 1659 1946 1663
rect 1958 1658 1962 1662
rect 1890 1650 1894 1654
rect 1890 1641 1894 1645
rect 1942 1651 1946 1655
rect 1958 1650 1962 1654
rect 1942 1642 1946 1646
rect 1958 1641 1962 1645
rect 1890 1633 1894 1637
rect 1942 1634 1946 1638
rect 1958 1633 1962 1637
rect 1890 1625 1894 1629
rect 1890 1616 1894 1620
rect 1942 1626 1946 1630
rect 1958 1625 1962 1629
rect 1942 1617 1946 1621
rect 1958 1616 1962 1620
rect 1890 1608 1894 1612
rect 1942 1609 1946 1613
rect 1958 1608 1962 1612
rect 1890 1600 1894 1604
rect 1890 1591 1894 1595
rect 1942 1601 1946 1605
rect 1958 1600 1962 1604
rect 1942 1592 1946 1596
rect 1958 1591 1962 1595
rect 1890 1583 1894 1587
rect 1942 1584 1946 1588
rect 1958 1583 1962 1587
rect 1890 1575 1894 1579
rect 1890 1566 1894 1570
rect 1942 1576 1946 1580
rect 1958 1575 1962 1579
rect 1942 1567 1946 1571
rect 1958 1566 1962 1570
rect 1890 1558 1894 1562
rect 1942 1559 1946 1563
rect 1958 1558 1962 1562
rect 1890 1550 1894 1554
rect 1890 1541 1894 1545
rect 1942 1551 1946 1555
rect 1958 1550 1962 1554
rect 1942 1542 1946 1546
rect 1958 1541 1962 1545
rect 1890 1533 1894 1537
rect 1942 1534 1946 1538
rect 1958 1533 1962 1537
rect 1890 1525 1894 1529
rect 1890 1516 1894 1520
rect 1942 1526 1946 1530
rect 1958 1525 1962 1529
rect 1942 1517 1946 1521
rect 1958 1516 1962 1520
rect 1890 1508 1894 1512
rect 1942 1509 1946 1513
rect 1958 1508 1962 1512
rect 1890 1500 1894 1504
rect 1890 1491 1894 1495
rect 1942 1501 1946 1505
rect 1958 1500 1962 1504
rect 1942 1492 1946 1496
rect 1958 1491 1962 1495
rect 1890 1483 1894 1487
rect 1942 1484 1946 1488
rect 1958 1483 1962 1487
rect 1890 1475 1894 1479
rect 1890 1466 1894 1470
rect 1942 1476 1946 1480
rect 1958 1475 1962 1479
rect 1942 1467 1946 1471
rect 1958 1466 1962 1470
rect 1890 1458 1894 1462
rect 1942 1459 1946 1463
rect 1958 1458 1962 1462
rect 1890 1450 1894 1454
rect 1890 1441 1894 1445
rect 1942 1451 1946 1455
rect 1958 1450 1962 1454
rect 1942 1442 1946 1446
rect 1958 1441 1962 1445
rect 1890 1433 1894 1437
rect 1942 1434 1946 1438
rect 1958 1433 1962 1437
rect 1890 1425 1894 1429
rect 1890 1416 1894 1420
rect 1942 1426 1946 1430
rect 1958 1425 1962 1429
rect 1942 1417 1946 1421
rect 1958 1416 1962 1420
rect 1890 1408 1894 1412
rect 1942 1409 1946 1413
rect 1958 1408 1962 1412
rect 1890 1400 1894 1404
rect 1890 1391 1894 1395
rect 1942 1401 1946 1405
rect 1958 1400 1962 1404
rect 1942 1392 1946 1396
rect 1958 1391 1962 1395
rect 1890 1383 1894 1387
rect 1942 1384 1946 1388
rect 1958 1383 1962 1387
rect 1752 1370 1756 1380
rect 1762 1370 1766 1380
rect 1890 1375 1894 1379
rect 1890 1366 1894 1370
rect 1942 1376 1946 1380
rect 1958 1375 1962 1379
rect 1942 1367 1946 1371
rect 1958 1366 1962 1370
rect 1890 1358 1894 1362
rect 1942 1359 1946 1363
rect 1958 1358 1962 1362
rect 1890 1350 1894 1354
rect 1890 1341 1894 1345
rect 1942 1351 1946 1355
rect 1958 1350 1962 1354
rect 1942 1342 1946 1346
rect 1958 1341 1962 1345
rect 1890 1333 1894 1337
rect 1942 1334 1946 1338
rect 1958 1333 1962 1337
rect 1890 1325 1894 1329
rect 1890 1316 1894 1320
rect 1942 1326 1946 1330
rect 1958 1325 1962 1329
rect 1942 1317 1946 1321
rect 1958 1316 1962 1320
rect 1890 1308 1894 1312
rect 1942 1309 1946 1313
rect 1958 1308 1962 1312
rect 1890 1300 1894 1304
rect 1890 1291 1894 1295
rect 1942 1301 1946 1305
rect 1958 1300 1962 1304
rect 1942 1292 1946 1296
rect 1958 1291 1962 1295
rect 1890 1283 1894 1287
rect 1942 1284 1946 1288
rect 1958 1283 1962 1287
rect 1890 1275 1894 1279
rect 1890 1266 1894 1270
rect 1942 1276 1946 1280
rect 1958 1275 1962 1279
rect 1942 1267 1946 1271
rect 1958 1266 1962 1270
rect 1890 1258 1894 1262
rect 1942 1259 1946 1263
rect 1958 1258 1962 1262
rect 1890 1250 1894 1254
rect 1890 1241 1894 1245
rect 1942 1251 1946 1255
rect 1958 1250 1962 1254
rect 1942 1242 1946 1246
rect 1958 1241 1962 1245
rect 1890 1233 1894 1237
rect 1942 1234 1946 1238
rect 1958 1233 1962 1237
rect 1890 1225 1894 1229
rect 1890 1216 1894 1220
rect 1942 1226 1946 1230
rect 1958 1225 1962 1229
rect 1942 1217 1946 1221
rect 1958 1216 1962 1220
rect 1890 1208 1894 1212
rect 1942 1209 1946 1213
rect 1958 1208 1962 1212
rect 1890 1200 1894 1204
rect 906 1188 910 1198
rect 916 1188 920 1198
rect 1890 1191 1894 1195
rect 1942 1201 1946 1205
rect 1958 1200 1962 1204
rect 1942 1192 1946 1196
rect 1958 1191 1962 1195
rect 1890 1183 1894 1187
rect 1942 1184 1946 1188
rect 1958 1183 1962 1187
rect 1890 1175 1894 1179
rect 1890 1166 1894 1170
rect 1942 1176 1946 1180
rect 1958 1175 1962 1179
rect 1942 1167 1946 1171
rect 1958 1166 1962 1170
rect 1890 1158 1894 1162
rect 1942 1159 1946 1163
rect 1958 1158 1962 1162
rect 1890 1150 1894 1154
rect 1890 1141 1894 1145
rect 1942 1151 1946 1155
rect 1958 1150 1962 1154
rect 1942 1142 1946 1146
rect 1958 1141 1962 1145
rect 1890 1133 1894 1137
rect 1942 1134 1946 1138
rect 1958 1133 1962 1137
rect 1890 1125 1894 1129
rect 1890 1116 1894 1120
rect 1942 1126 1946 1130
rect 1958 1125 1962 1129
rect 1942 1117 1946 1121
rect 1958 1116 1962 1120
rect 1890 1108 1894 1112
rect 1942 1109 1946 1113
rect 1958 1108 1962 1112
rect 1890 1100 1894 1104
rect 1890 1091 1894 1095
rect 1942 1101 1946 1105
rect 1958 1100 1962 1104
rect 1942 1092 1946 1096
rect 1958 1091 1962 1095
rect 1890 1083 1894 1087
rect 1942 1084 1946 1088
rect 1958 1083 1962 1087
rect 1890 1075 1894 1079
rect 1890 1066 1894 1070
rect 1942 1076 1946 1080
rect 1958 1075 1962 1079
rect 1942 1067 1946 1071
rect 1958 1066 1962 1070
rect 1729 1055 1733 1065
rect 1739 1055 1743 1065
rect 1747 1055 1751 1065
rect 1757 1055 1761 1065
rect 1767 1055 1771 1065
rect 1890 1058 1894 1062
rect 1942 1059 1946 1063
rect 1958 1058 1962 1062
rect 1890 1050 1894 1054
rect 1890 1041 1894 1045
rect 1942 1051 1946 1055
rect 1958 1050 1962 1054
rect 1942 1042 1946 1046
rect 1958 1041 1962 1045
rect 1890 1033 1894 1037
rect 1942 1034 1946 1038
rect 1958 1033 1962 1037
rect 1890 1025 1894 1029
rect 1890 1016 1894 1020
rect 1942 1026 1946 1030
rect 1958 1025 1962 1029
rect 1942 1017 1946 1021
rect 1958 1016 1962 1020
rect 1890 1008 1894 1012
rect 1942 1009 1946 1013
rect 1958 1008 1962 1012
rect 1890 1000 1894 1004
rect 1890 991 1894 995
rect 1942 1001 1946 1005
rect 1958 1000 1962 1004
rect 1942 992 1946 996
rect 1958 991 1962 995
rect 1890 983 1894 987
rect 1942 984 1946 988
rect 1958 983 1962 987
rect 1890 975 1894 979
rect 1890 966 1894 970
rect 1942 976 1946 980
rect 1958 975 1962 979
rect 1942 967 1946 971
rect 1958 966 1962 970
rect 1890 958 1894 962
rect 1942 959 1946 963
rect 1958 958 1962 962
rect 1890 950 1894 954
rect 1890 941 1894 945
rect 1942 951 1946 955
rect 1958 950 1962 954
rect 1942 942 1946 946
rect 1958 941 1962 945
rect 1890 933 1894 937
rect 1942 934 1946 938
rect 1958 933 1962 937
rect 1890 925 1894 929
rect 1890 916 1894 920
rect 1942 926 1946 930
rect 1958 925 1962 929
rect 1942 917 1946 921
rect 1958 916 1962 920
rect 1890 908 1894 912
rect 1942 909 1946 913
rect 1958 908 1962 912
rect 1890 900 1894 904
rect 1890 891 1894 895
rect 1942 901 1946 905
rect 1958 900 1962 904
rect 1942 892 1946 896
rect 1958 891 1962 895
rect 1890 883 1894 887
rect 1942 884 1946 888
rect 1958 883 1962 887
rect 1890 875 1894 879
rect 1890 866 1894 870
rect 1942 876 1946 880
rect 1958 875 1962 879
rect 1942 867 1946 871
rect 1958 866 1962 870
rect 1890 858 1894 862
rect 1942 859 1946 863
rect 1958 858 1962 862
rect 1890 850 1894 854
rect 1890 841 1894 845
rect 1942 851 1946 855
rect 1958 850 1962 854
rect 1942 842 1946 846
rect 1958 841 1962 845
rect 1890 833 1894 837
rect 1942 834 1946 838
rect 1958 833 1962 837
rect 1890 825 1894 829
rect 1890 816 1894 820
rect 1942 826 1946 830
rect 1958 825 1962 829
rect 1942 817 1946 821
rect 1958 816 1962 820
rect 1890 808 1894 812
rect 1942 809 1946 813
rect 1958 808 1962 812
rect 1890 800 1894 804
rect 1890 791 1894 795
rect 1942 801 1946 805
rect 1958 800 1962 804
rect 1942 792 1946 796
rect 1958 791 1962 795
rect 1890 783 1894 787
rect 1942 784 1946 788
rect 1958 783 1962 787
rect 1890 775 1894 779
rect 1890 766 1894 770
rect 1942 776 1946 780
rect 1958 775 1962 779
rect 1942 767 1946 771
rect 1958 766 1962 770
rect 1890 758 1894 762
rect 1942 759 1946 763
rect 1958 758 1962 762
rect 1890 750 1894 754
rect 1890 741 1894 745
rect 1942 751 1946 755
rect 1958 750 1962 754
rect 1942 742 1946 746
rect 1958 741 1962 745
rect 1890 733 1894 737
rect 1942 734 1946 738
rect 1958 733 1962 737
rect 1890 725 1894 729
rect 1890 716 1894 720
rect 1942 726 1946 730
rect 1958 725 1962 729
rect 1942 717 1946 721
rect 1958 716 1962 720
rect 1890 708 1894 712
rect 1942 709 1946 713
rect 1958 708 1962 712
rect 1890 700 1894 704
rect 1890 691 1894 695
rect 1942 701 1946 705
rect 1958 700 1962 704
rect 1942 692 1946 696
rect 1958 691 1962 695
rect 1890 683 1894 687
rect 1942 684 1946 688
rect 1958 683 1962 687
rect 1890 675 1894 679
rect 1890 666 1894 670
rect 1942 676 1946 680
rect 1958 675 1962 679
rect 1942 667 1946 671
rect 1958 666 1962 670
rect 1890 658 1894 662
rect 1942 659 1946 663
rect 1958 658 1962 662
rect 1890 650 1894 654
rect 1890 641 1894 645
rect 1942 651 1946 655
rect 1958 650 1962 654
rect 1942 642 1946 646
rect 1958 641 1962 645
rect 1890 633 1894 637
rect 1942 634 1946 638
rect 1958 633 1962 637
rect 1890 625 1894 629
rect 1890 616 1894 620
rect 1942 626 1946 630
rect 1958 625 1962 629
rect 1942 617 1946 621
rect 1958 616 1962 620
rect 1890 608 1894 612
rect 1942 609 1946 613
rect 1958 608 1962 612
rect 1890 600 1894 604
rect 1890 591 1894 595
rect 1942 601 1946 605
rect 1958 600 1962 604
rect 1942 592 1946 596
rect 1958 591 1962 595
rect 1890 583 1894 587
rect 1942 584 1946 588
rect 1958 583 1962 587
rect 1890 575 1894 579
rect 1890 566 1894 570
rect 1942 576 1946 580
rect 1958 575 1962 579
rect 1942 567 1946 571
rect 1958 566 1962 570
rect 1890 558 1894 562
rect 1942 559 1946 563
rect 1958 558 1962 562
rect 1890 550 1894 554
rect 1890 541 1894 545
rect 1942 551 1946 555
rect 1958 550 1962 554
rect 1942 542 1946 546
rect 1958 541 1962 545
rect 1890 533 1894 537
rect 1942 534 1946 538
rect 1958 533 1962 537
rect 1890 525 1894 529
rect 1890 516 1894 520
rect 1942 526 1946 530
rect 1958 525 1962 529
rect 1942 517 1946 521
rect 1958 516 1962 520
rect 1890 508 1894 512
rect 1942 509 1946 513
rect 1958 508 1962 512
rect 1890 500 1894 504
rect 1890 491 1894 495
rect 1942 501 1946 505
rect 1958 500 1962 504
rect 1942 492 1946 496
rect 1958 491 1962 495
rect 1890 483 1894 487
rect 1942 484 1946 488
rect 1958 483 1962 487
rect 1890 475 1894 479
rect 1890 466 1894 470
rect 1942 476 1946 480
rect 1958 475 1962 479
rect 1942 467 1946 471
rect 1958 466 1962 470
rect 1890 458 1894 462
rect 1942 459 1946 463
rect 1958 458 1962 462
rect 1890 450 1894 454
rect 1890 441 1894 445
rect 1942 451 1946 455
rect 1958 450 1962 454
rect 1942 442 1946 446
rect 1958 441 1962 445
rect 1890 433 1894 437
rect 1942 434 1946 438
rect 1958 433 1962 437
rect 1890 425 1894 429
rect 1890 416 1894 420
rect 1942 426 1946 430
rect 1958 425 1962 429
rect 1942 417 1946 421
rect 1958 416 1962 420
rect 1890 408 1894 412
rect 1942 409 1946 413
rect 1958 408 1962 412
rect 1890 400 1894 404
rect 1890 391 1894 395
rect 1942 401 1946 405
rect 1958 400 1962 404
rect 1942 392 1946 396
rect 1958 391 1962 395
rect 1890 383 1894 387
rect 1942 384 1946 388
rect 1958 383 1962 387
rect 1890 375 1894 379
rect 1890 366 1894 370
rect 1942 376 1946 380
rect 1958 375 1962 379
rect 1942 367 1946 371
rect 1958 366 1962 370
rect 1890 358 1894 362
rect 1942 359 1946 363
rect 1958 358 1962 362
rect 1890 350 1894 354
rect 1890 341 1894 345
rect 1942 351 1946 355
rect 1958 350 1962 354
rect 1942 342 1946 346
rect 1958 341 1962 345
rect 1890 333 1894 337
rect 1942 334 1946 338
rect 1958 333 1962 337
rect 1890 325 1894 329
rect 1890 316 1894 320
rect 1942 326 1946 330
rect 1958 325 1962 329
rect 1942 317 1946 321
rect 1958 316 1962 320
rect 1890 308 1894 312
rect 1942 309 1946 313
rect 1958 308 1962 312
rect 1890 300 1894 304
rect 1890 291 1894 295
rect 1942 301 1946 305
rect 1958 300 1962 304
rect 1942 292 1946 296
rect 1958 291 1962 295
rect 1890 283 1894 287
rect 1942 284 1946 288
rect 1958 283 1962 287
rect 1890 275 1894 279
rect 1890 266 1894 270
rect 1942 276 1946 280
rect 1958 275 1962 279
rect 1942 267 1946 271
rect 1958 266 1962 270
rect 1890 258 1894 262
rect 1942 259 1946 263
rect 1958 258 1962 262
rect 1890 250 1894 254
rect 1890 241 1894 245
rect 1942 251 1946 255
rect 1958 250 1962 254
rect 1942 242 1946 246
rect 1958 241 1962 245
rect 1890 233 1894 237
rect 1942 234 1946 238
rect 1958 233 1962 237
rect 1890 225 1894 229
rect 1890 216 1894 220
rect 1942 226 1946 230
rect 1958 225 1962 229
rect 1942 217 1946 221
rect 1958 216 1962 220
rect 1890 208 1894 212
rect 1942 209 1946 213
rect 1958 208 1962 212
rect 1890 200 1894 204
rect 1890 191 1894 195
rect 1942 201 1946 205
rect 1958 200 1962 204
rect 1942 192 1946 196
rect 1958 191 1962 195
rect 1890 183 1894 187
rect 1942 184 1946 188
rect 1958 183 1962 187
rect 1890 175 1894 179
rect 1890 166 1894 170
rect 1942 176 1946 180
rect 1958 175 1962 179
rect 1942 167 1946 171
rect 1958 166 1962 170
rect 1890 158 1894 162
rect 1942 159 1946 163
rect 1958 158 1962 162
rect 1890 150 1894 154
rect 1890 141 1894 145
rect 1942 151 1946 155
rect 1958 150 1962 154
rect 1942 142 1946 146
rect 1958 141 1962 145
rect 1890 133 1894 137
rect 1942 134 1946 138
rect 1958 133 1962 137
rect 1890 125 1894 129
rect 1890 116 1894 120
rect 1942 126 1946 130
rect 1958 125 1962 129
rect 1942 117 1946 121
rect 1958 116 1962 120
rect 1890 108 1894 112
rect 1942 109 1946 113
rect 1958 108 1962 112
rect 1890 100 1894 104
rect 1890 91 1894 95
rect 1942 101 1946 105
rect 1958 100 1962 104
rect 1942 92 1946 96
rect 1958 91 1962 95
rect 1890 83 1894 87
rect 1942 84 1946 88
rect 1958 83 1962 87
rect 1890 75 1894 79
rect 1890 66 1894 70
rect 1942 76 1946 80
rect 1958 75 1962 79
rect 1942 67 1946 71
rect 1958 66 1962 70
rect 1890 58 1894 62
rect 1942 59 1946 63
rect 1958 58 1962 62
rect 1890 50 1894 54
rect 1890 41 1894 45
rect 1942 51 1946 55
rect 1958 50 1962 54
rect 1942 42 1946 46
rect 1958 41 1962 45
rect 1890 33 1894 37
rect 1942 34 1946 38
rect 1958 33 1962 37
rect 1890 25 1894 29
rect 1942 26 1946 30
rect 1958 25 1962 29
<< pdcontact >>
rect 1904 2016 1912 2020
rect 1924 2017 1932 2021
rect 1904 2008 1912 2012
rect 1924 2009 1932 2013
rect 1972 2016 1980 2020
rect 1904 2000 1912 2004
rect 1924 2001 1932 2005
rect 1972 2008 1980 2012
rect 1904 1991 1912 1995
rect 1924 1992 1932 1996
rect 1972 2000 1980 2004
rect 1904 1983 1912 1987
rect 1924 1984 1932 1988
rect 1972 1991 1980 1995
rect 1904 1975 1912 1979
rect 1924 1976 1932 1980
rect 1972 1983 1980 1987
rect 1904 1966 1912 1970
rect 1924 1967 1932 1971
rect 1972 1975 1980 1979
rect 1904 1958 1912 1962
rect 1924 1959 1932 1963
rect 1972 1966 1980 1970
rect 1904 1950 1912 1954
rect 1924 1951 1932 1955
rect 1972 1958 1980 1962
rect 1904 1941 1912 1945
rect 1924 1942 1932 1946
rect 1972 1950 1980 1954
rect 1904 1933 1912 1937
rect 1924 1934 1932 1938
rect 1972 1941 1980 1945
rect 1904 1925 1912 1929
rect 1924 1926 1932 1930
rect 1972 1933 1980 1937
rect 1904 1916 1912 1920
rect 1924 1917 1932 1921
rect 1972 1925 1980 1929
rect 1904 1908 1912 1912
rect 1924 1909 1932 1913
rect 1972 1916 1980 1920
rect 1904 1900 1912 1904
rect 1924 1901 1932 1905
rect 1972 1908 1980 1912
rect 1904 1891 1912 1895
rect 1924 1892 1932 1896
rect 1972 1900 1980 1904
rect 1904 1883 1912 1887
rect 1924 1884 1932 1888
rect 1972 1891 1980 1895
rect 1904 1875 1912 1879
rect 1924 1876 1932 1880
rect 1972 1883 1980 1887
rect 1904 1866 1912 1870
rect 1924 1867 1932 1871
rect 1972 1875 1980 1879
rect 1904 1858 1912 1862
rect 1924 1859 1932 1863
rect 1972 1866 1980 1870
rect 1904 1850 1912 1854
rect 1924 1851 1932 1855
rect 1972 1858 1980 1862
rect 1904 1841 1912 1845
rect 1924 1842 1932 1846
rect 1972 1850 1980 1854
rect 1904 1833 1912 1837
rect 1924 1834 1932 1838
rect 1972 1841 1980 1845
rect 1904 1825 1912 1829
rect 1924 1826 1932 1830
rect 1972 1833 1980 1837
rect 1904 1816 1912 1820
rect 1924 1817 1932 1821
rect 1972 1825 1980 1829
rect 1904 1808 1912 1812
rect 1924 1809 1932 1813
rect 1972 1816 1980 1820
rect 1904 1800 1912 1804
rect 1924 1801 1932 1805
rect 1972 1808 1980 1812
rect 1904 1791 1912 1795
rect 1924 1792 1932 1796
rect 1972 1800 1980 1804
rect 1904 1783 1912 1787
rect 1924 1784 1932 1788
rect 1972 1791 1980 1795
rect 1904 1775 1912 1779
rect 1924 1776 1932 1780
rect 1972 1783 1980 1787
rect 1904 1766 1912 1770
rect 1924 1767 1932 1771
rect 1972 1775 1980 1779
rect 1904 1758 1912 1762
rect 1924 1759 1932 1763
rect 1972 1766 1980 1770
rect 1904 1750 1912 1754
rect 1924 1751 1932 1755
rect 1972 1758 1980 1762
rect 1904 1741 1912 1745
rect 1924 1742 1932 1746
rect 1972 1750 1980 1754
rect 1904 1733 1912 1737
rect 1924 1734 1932 1738
rect 1972 1741 1980 1745
rect 1904 1725 1912 1729
rect 1924 1726 1932 1730
rect 1972 1733 1980 1737
rect 1904 1716 1912 1720
rect 1924 1717 1932 1721
rect 1972 1725 1980 1729
rect 1904 1708 1912 1712
rect 1924 1709 1932 1713
rect 1972 1716 1980 1720
rect 1904 1700 1912 1704
rect 1924 1701 1932 1705
rect 1972 1708 1980 1712
rect 1904 1691 1912 1695
rect 1924 1692 1932 1696
rect 1972 1700 1980 1704
rect 1904 1683 1912 1687
rect 1924 1684 1932 1688
rect 1972 1691 1980 1695
rect 1904 1675 1912 1679
rect 1924 1676 1932 1680
rect 1972 1683 1980 1687
rect 1904 1666 1912 1670
rect 1924 1667 1932 1671
rect 1972 1675 1980 1679
rect 1904 1658 1912 1662
rect 1924 1659 1932 1663
rect 1972 1666 1980 1670
rect 1904 1650 1912 1654
rect 1924 1651 1932 1655
rect 1972 1658 1980 1662
rect 1904 1641 1912 1645
rect 1924 1642 1932 1646
rect 1972 1650 1980 1654
rect 1904 1633 1912 1637
rect 1924 1634 1932 1638
rect 1972 1641 1980 1645
rect 1904 1625 1912 1629
rect 1924 1626 1932 1630
rect 1972 1633 1980 1637
rect 1904 1616 1912 1620
rect 1924 1617 1932 1621
rect 1972 1625 1980 1629
rect 1904 1608 1912 1612
rect 1924 1609 1932 1613
rect 1972 1616 1980 1620
rect 1904 1600 1912 1604
rect 1924 1601 1932 1605
rect 1972 1608 1980 1612
rect 1904 1591 1912 1595
rect 1924 1592 1932 1596
rect 1972 1600 1980 1604
rect 1904 1583 1912 1587
rect 1924 1584 1932 1588
rect 1972 1591 1980 1595
rect 1904 1575 1912 1579
rect 1924 1576 1932 1580
rect 1972 1583 1980 1587
rect 1904 1566 1912 1570
rect 1924 1567 1932 1571
rect 1972 1575 1980 1579
rect 1904 1558 1912 1562
rect 1924 1559 1932 1563
rect 1972 1566 1980 1570
rect 1904 1550 1912 1554
rect 1924 1551 1932 1555
rect 1972 1558 1980 1562
rect 1904 1541 1912 1545
rect 1924 1542 1932 1546
rect 1972 1550 1980 1554
rect 1904 1533 1912 1537
rect 1924 1534 1932 1538
rect 1972 1541 1980 1545
rect 1904 1525 1912 1529
rect 1924 1526 1932 1530
rect 1972 1533 1980 1537
rect 1904 1516 1912 1520
rect 1924 1517 1932 1521
rect 1972 1525 1980 1529
rect 1904 1508 1912 1512
rect 1924 1509 1932 1513
rect 1972 1516 1980 1520
rect 1904 1500 1912 1504
rect 1924 1501 1932 1505
rect 1972 1508 1980 1512
rect 1904 1491 1912 1495
rect 1924 1492 1932 1496
rect 1972 1500 1980 1504
rect 1904 1483 1912 1487
rect 1924 1484 1932 1488
rect 1972 1491 1980 1495
rect 1904 1475 1912 1479
rect 1924 1476 1932 1480
rect 1972 1483 1980 1487
rect 1904 1466 1912 1470
rect 1924 1467 1932 1471
rect 1972 1475 1980 1479
rect 1904 1458 1912 1462
rect 1924 1459 1932 1463
rect 1972 1466 1980 1470
rect 1904 1450 1912 1454
rect 1924 1451 1932 1455
rect 1972 1458 1980 1462
rect 1904 1441 1912 1445
rect 1924 1442 1932 1446
rect 1972 1450 1980 1454
rect 1904 1433 1912 1437
rect 1924 1434 1932 1438
rect 1972 1441 1980 1445
rect 1904 1425 1912 1429
rect 1924 1426 1932 1430
rect 1972 1433 1980 1437
rect 1904 1416 1912 1420
rect 1924 1417 1932 1421
rect 1972 1425 1980 1429
rect 1752 1390 1756 1410
rect 1762 1390 1766 1410
rect 1904 1408 1912 1412
rect 1924 1409 1932 1413
rect 1972 1416 1980 1420
rect 1904 1400 1912 1404
rect 1924 1401 1932 1405
rect 1972 1408 1980 1412
rect 1904 1391 1912 1395
rect 1924 1392 1932 1396
rect 1972 1400 1980 1404
rect 1904 1383 1912 1387
rect 1924 1384 1932 1388
rect 1972 1391 1980 1395
rect 1904 1375 1912 1379
rect 1924 1376 1932 1380
rect 1972 1383 1980 1387
rect 1904 1366 1912 1370
rect 1924 1367 1932 1371
rect 1972 1375 1980 1379
rect 1904 1358 1912 1362
rect 1924 1359 1932 1363
rect 1972 1366 1980 1370
rect 1904 1350 1912 1354
rect 1924 1351 1932 1355
rect 1972 1358 1980 1362
rect 1904 1341 1912 1345
rect 1924 1342 1932 1346
rect 1972 1350 1980 1354
rect 1904 1333 1912 1337
rect 1924 1334 1932 1338
rect 1972 1341 1980 1345
rect 1904 1325 1912 1329
rect 1924 1326 1932 1330
rect 1972 1333 1980 1337
rect 1904 1316 1912 1320
rect 1924 1317 1932 1321
rect 1972 1325 1980 1329
rect 1904 1308 1912 1312
rect 1924 1309 1932 1313
rect 1972 1316 1980 1320
rect 1904 1300 1912 1304
rect 1924 1301 1932 1305
rect 1972 1308 1980 1312
rect 1904 1291 1912 1295
rect 1924 1292 1932 1296
rect 1972 1300 1980 1304
rect 1904 1283 1912 1287
rect 1924 1284 1932 1288
rect 1972 1291 1980 1295
rect 1904 1275 1912 1279
rect 1924 1276 1932 1280
rect 1972 1283 1980 1287
rect 1904 1266 1912 1270
rect 1924 1267 1932 1271
rect 1972 1275 1980 1279
rect 1904 1258 1912 1262
rect 1924 1259 1932 1263
rect 1972 1266 1980 1270
rect 1904 1250 1912 1254
rect 1924 1251 1932 1255
rect 1972 1258 1980 1262
rect 1904 1241 1912 1245
rect 1924 1242 1932 1246
rect 1972 1250 1980 1254
rect 1904 1233 1912 1237
rect 1924 1234 1932 1238
rect 1972 1241 1980 1245
rect 1904 1225 1912 1229
rect 1924 1226 1932 1230
rect 1972 1233 1980 1237
rect 1904 1216 1912 1220
rect 1924 1217 1932 1221
rect 1972 1225 1980 1229
rect 1904 1208 1912 1212
rect 1924 1209 1932 1213
rect 1972 1216 1980 1220
rect 1904 1200 1912 1204
rect 1924 1201 1932 1205
rect 1972 1208 1980 1212
rect 1904 1191 1912 1195
rect 1924 1192 1932 1196
rect 1972 1200 1980 1204
rect 1904 1183 1912 1187
rect 1924 1184 1932 1188
rect 1972 1191 1980 1195
rect 906 1158 910 1178
rect 916 1158 920 1178
rect 1904 1175 1912 1179
rect 1924 1176 1932 1180
rect 1972 1183 1980 1187
rect 1904 1166 1912 1170
rect 1924 1167 1932 1171
rect 1972 1175 1980 1179
rect 1904 1158 1912 1162
rect 1924 1159 1932 1163
rect 1972 1166 1980 1170
rect 1904 1150 1912 1154
rect 1924 1151 1932 1155
rect 1972 1158 1980 1162
rect 1904 1141 1912 1145
rect 1924 1142 1932 1146
rect 1972 1150 1980 1154
rect 1904 1133 1912 1137
rect 1924 1134 1932 1138
rect 1972 1141 1980 1145
rect 1904 1125 1912 1129
rect 1924 1126 1932 1130
rect 1972 1133 1980 1137
rect 1904 1116 1912 1120
rect 1924 1117 1932 1121
rect 1972 1125 1980 1129
rect 1904 1108 1912 1112
rect 1924 1109 1932 1113
rect 1972 1116 1980 1120
rect 1904 1100 1912 1104
rect 1924 1101 1932 1105
rect 1729 1075 1733 1093
rect 1739 1075 1743 1093
rect 1747 1075 1751 1093
rect 1757 1075 1761 1093
rect 1767 1075 1771 1093
rect 1972 1108 1980 1112
rect 1904 1091 1912 1095
rect 1924 1092 1932 1096
rect 1972 1100 1980 1104
rect 1904 1083 1912 1087
rect 1924 1084 1932 1088
rect 1972 1091 1980 1095
rect 1904 1075 1912 1079
rect 1924 1076 1932 1080
rect 1972 1083 1980 1087
rect 1904 1066 1912 1070
rect 1924 1067 1932 1071
rect 1972 1075 1980 1079
rect 1904 1058 1912 1062
rect 1924 1059 1932 1063
rect 1972 1066 1980 1070
rect 1904 1050 1912 1054
rect 1924 1051 1932 1055
rect 1972 1058 1980 1062
rect 1904 1041 1912 1045
rect 1924 1042 1932 1046
rect 1972 1050 1980 1054
rect 1904 1033 1912 1037
rect 1924 1034 1932 1038
rect 1972 1041 1980 1045
rect 1904 1025 1912 1029
rect 1924 1026 1932 1030
rect 1972 1033 1980 1037
rect 1904 1016 1912 1020
rect 1924 1017 1932 1021
rect 1972 1025 1980 1029
rect 1904 1008 1912 1012
rect 1924 1009 1932 1013
rect 1972 1016 1980 1020
rect 1904 1000 1912 1004
rect 1924 1001 1932 1005
rect 1972 1008 1980 1012
rect 1904 991 1912 995
rect 1924 992 1932 996
rect 1972 1000 1980 1004
rect 1904 983 1912 987
rect 1924 984 1932 988
rect 1972 991 1980 995
rect 1904 975 1912 979
rect 1924 976 1932 980
rect 1972 983 1980 987
rect 1904 966 1912 970
rect 1924 967 1932 971
rect 1972 975 1980 979
rect 1904 958 1912 962
rect 1924 959 1932 963
rect 1972 966 1980 970
rect 1904 950 1912 954
rect 1924 951 1932 955
rect 1972 958 1980 962
rect 1904 941 1912 945
rect 1924 942 1932 946
rect 1972 950 1980 954
rect 1904 933 1912 937
rect 1924 934 1932 938
rect 1972 941 1980 945
rect 1904 925 1912 929
rect 1924 926 1932 930
rect 1972 933 1980 937
rect 1904 916 1912 920
rect 1924 917 1932 921
rect 1972 925 1980 929
rect 1904 908 1912 912
rect 1924 909 1932 913
rect 1972 916 1980 920
rect 1904 900 1912 904
rect 1924 901 1932 905
rect 1972 908 1980 912
rect 1904 891 1912 895
rect 1924 892 1932 896
rect 1972 900 1980 904
rect 1904 883 1912 887
rect 1924 884 1932 888
rect 1972 891 1980 895
rect 1904 875 1912 879
rect 1924 876 1932 880
rect 1972 883 1980 887
rect 1904 866 1912 870
rect 1924 867 1932 871
rect 1972 875 1980 879
rect 1904 858 1912 862
rect 1924 859 1932 863
rect 1972 866 1980 870
rect 1904 850 1912 854
rect 1924 851 1932 855
rect 1972 858 1980 862
rect 1904 841 1912 845
rect 1924 842 1932 846
rect 1972 850 1980 854
rect 1904 833 1912 837
rect 1924 834 1932 838
rect 1972 841 1980 845
rect 1904 825 1912 829
rect 1924 826 1932 830
rect 1972 833 1980 837
rect 1904 816 1912 820
rect 1924 817 1932 821
rect 1972 825 1980 829
rect 1904 808 1912 812
rect 1924 809 1932 813
rect 1972 816 1980 820
rect 1904 800 1912 804
rect 1924 801 1932 805
rect 1972 808 1980 812
rect 1904 791 1912 795
rect 1924 792 1932 796
rect 1972 800 1980 804
rect 1904 783 1912 787
rect 1924 784 1932 788
rect 1972 791 1980 795
rect 1904 775 1912 779
rect 1924 776 1932 780
rect 1972 783 1980 787
rect 1904 766 1912 770
rect 1924 767 1932 771
rect 1972 775 1980 779
rect 1904 758 1912 762
rect 1924 759 1932 763
rect 1972 766 1980 770
rect 1904 750 1912 754
rect 1924 751 1932 755
rect 1972 758 1980 762
rect 1904 741 1912 745
rect 1924 742 1932 746
rect 1972 750 1980 754
rect 1904 733 1912 737
rect 1924 734 1932 738
rect 1972 741 1980 745
rect 1904 725 1912 729
rect 1924 726 1932 730
rect 1972 733 1980 737
rect 1904 716 1912 720
rect 1924 717 1932 721
rect 1972 725 1980 729
rect 1904 708 1912 712
rect 1924 709 1932 713
rect 1972 716 1980 720
rect 1904 700 1912 704
rect 1924 701 1932 705
rect 1972 708 1980 712
rect 1904 691 1912 695
rect 1924 692 1932 696
rect 1972 700 1980 704
rect 1904 683 1912 687
rect 1924 684 1932 688
rect 1972 691 1980 695
rect 1904 675 1912 679
rect 1924 676 1932 680
rect 1972 683 1980 687
rect 1904 666 1912 670
rect 1924 667 1932 671
rect 1972 675 1980 679
rect 1904 658 1912 662
rect 1924 659 1932 663
rect 1972 666 1980 670
rect 1904 650 1912 654
rect 1924 651 1932 655
rect 1972 658 1980 662
rect 1904 641 1912 645
rect 1924 642 1932 646
rect 1972 650 1980 654
rect 1904 633 1912 637
rect 1924 634 1932 638
rect 1972 641 1980 645
rect 1904 625 1912 629
rect 1924 626 1932 630
rect 1972 633 1980 637
rect 1904 616 1912 620
rect 1924 617 1932 621
rect 1972 625 1980 629
rect 1904 608 1912 612
rect 1924 609 1932 613
rect 1972 616 1980 620
rect 1904 600 1912 604
rect 1924 601 1932 605
rect 1972 608 1980 612
rect 1904 591 1912 595
rect 1924 592 1932 596
rect 1972 600 1980 604
rect 1904 583 1912 587
rect 1924 584 1932 588
rect 1972 591 1980 595
rect 1904 575 1912 579
rect 1924 576 1932 580
rect 1972 583 1980 587
rect 1904 566 1912 570
rect 1924 567 1932 571
rect 1972 575 1980 579
rect 1904 558 1912 562
rect 1924 559 1932 563
rect 1972 566 1980 570
rect 1904 550 1912 554
rect 1924 551 1932 555
rect 1972 558 1980 562
rect 1904 541 1912 545
rect 1924 542 1932 546
rect 1972 550 1980 554
rect 1904 533 1912 537
rect 1924 534 1932 538
rect 1972 541 1980 545
rect 1904 525 1912 529
rect 1924 526 1932 530
rect 1972 533 1980 537
rect 1904 516 1912 520
rect 1924 517 1932 521
rect 1972 525 1980 529
rect 1904 508 1912 512
rect 1924 509 1932 513
rect 1972 516 1980 520
rect 1904 500 1912 504
rect 1924 501 1932 505
rect 1972 508 1980 512
rect 1904 491 1912 495
rect 1924 492 1932 496
rect 1972 500 1980 504
rect 1904 483 1912 487
rect 1924 484 1932 488
rect 1972 491 1980 495
rect 1904 475 1912 479
rect 1924 476 1932 480
rect 1972 483 1980 487
rect 1904 466 1912 470
rect 1924 467 1932 471
rect 1972 475 1980 479
rect 1904 458 1912 462
rect 1924 459 1932 463
rect 1972 466 1980 470
rect 1904 450 1912 454
rect 1924 451 1932 455
rect 1972 458 1980 462
rect 1904 441 1912 445
rect 1924 442 1932 446
rect 1972 450 1980 454
rect 1904 433 1912 437
rect 1924 434 1932 438
rect 1972 441 1980 445
rect 1904 425 1912 429
rect 1924 426 1932 430
rect 1972 433 1980 437
rect 1904 416 1912 420
rect 1924 417 1932 421
rect 1972 425 1980 429
rect 1904 408 1912 412
rect 1924 409 1932 413
rect 1972 416 1980 420
rect 1904 400 1912 404
rect 1924 401 1932 405
rect 1972 408 1980 412
rect 1904 391 1912 395
rect 1924 392 1932 396
rect 1972 400 1980 404
rect 1904 383 1912 387
rect 1924 384 1932 388
rect 1972 391 1980 395
rect 1904 375 1912 379
rect 1924 376 1932 380
rect 1972 383 1980 387
rect 1904 366 1912 370
rect 1924 367 1932 371
rect 1972 375 1980 379
rect 1904 358 1912 362
rect 1924 359 1932 363
rect 1972 366 1980 370
rect 1904 350 1912 354
rect 1924 351 1932 355
rect 1972 358 1980 362
rect 1904 341 1912 345
rect 1924 342 1932 346
rect 1972 350 1980 354
rect 1904 333 1912 337
rect 1924 334 1932 338
rect 1972 341 1980 345
rect 1904 325 1912 329
rect 1924 326 1932 330
rect 1972 333 1980 337
rect 1904 316 1912 320
rect 1924 317 1932 321
rect 1972 325 1980 329
rect 1904 308 1912 312
rect 1924 309 1932 313
rect 1972 316 1980 320
rect 1904 300 1912 304
rect 1924 301 1932 305
rect 1972 308 1980 312
rect 1904 291 1912 295
rect 1924 292 1932 296
rect 1972 300 1980 304
rect 1904 283 1912 287
rect 1924 284 1932 288
rect 1972 291 1980 295
rect 1904 275 1912 279
rect 1924 276 1932 280
rect 1972 283 1980 287
rect 1904 266 1912 270
rect 1924 267 1932 271
rect 1972 275 1980 279
rect 1904 258 1912 262
rect 1924 259 1932 263
rect 1972 266 1980 270
rect 1904 250 1912 254
rect 1924 251 1932 255
rect 1972 258 1980 262
rect 1904 241 1912 245
rect 1924 242 1932 246
rect 1972 250 1980 254
rect 1904 233 1912 237
rect 1924 234 1932 238
rect 1972 241 1980 245
rect 1904 225 1912 229
rect 1924 226 1932 230
rect 1972 233 1980 237
rect 1904 216 1912 220
rect 1924 217 1932 221
rect 1972 225 1980 229
rect 1904 208 1912 212
rect 1924 209 1932 213
rect 1972 216 1980 220
rect 1904 200 1912 204
rect 1924 201 1932 205
rect 1972 208 1980 212
rect 1904 191 1912 195
rect 1924 192 1932 196
rect 1972 200 1980 204
rect 1904 183 1912 187
rect 1924 184 1932 188
rect 1972 191 1980 195
rect 1904 175 1912 179
rect 1924 176 1932 180
rect 1972 183 1980 187
rect 1904 166 1912 170
rect 1924 167 1932 171
rect 1972 175 1980 179
rect 1904 158 1912 162
rect 1924 159 1932 163
rect 1972 166 1980 170
rect 1904 150 1912 154
rect 1924 151 1932 155
rect 1972 158 1980 162
rect 1904 141 1912 145
rect 1924 142 1932 146
rect 1972 150 1980 154
rect 1904 133 1912 137
rect 1924 134 1932 138
rect 1972 141 1980 145
rect 1904 125 1912 129
rect 1924 126 1932 130
rect 1972 133 1980 137
rect 1904 116 1912 120
rect 1924 117 1932 121
rect 1972 125 1980 129
rect 1904 108 1912 112
rect 1924 109 1932 113
rect 1972 116 1980 120
rect 1904 100 1912 104
rect 1924 101 1932 105
rect 1972 108 1980 112
rect 1904 91 1912 95
rect 1924 92 1932 96
rect 1972 100 1980 104
rect 1904 83 1912 87
rect 1924 84 1932 88
rect 1972 91 1980 95
rect 1904 75 1912 79
rect 1924 76 1932 80
rect 1972 83 1980 87
rect 1904 66 1912 70
rect 1924 67 1932 71
rect 1972 75 1980 79
rect 1904 58 1912 62
rect 1924 59 1932 63
rect 1972 66 1980 70
rect 1904 50 1912 54
rect 1924 51 1932 55
rect 1972 58 1980 62
rect 1904 41 1912 45
rect 1924 42 1932 46
rect 1972 50 1980 54
rect 1904 33 1912 37
rect 1924 34 1932 38
rect 1972 41 1980 45
rect 1904 25 1912 29
rect 1924 26 1932 30
rect 1972 33 1980 37
rect 1972 25 1980 29
<< m2contact >>
rect 920 2006 928 2014
rect 12 1880 20 1888
rect 43 1828 49 1833
rect 153 1829 159 1834
rect 263 1828 269 1833
rect 373 1829 379 1834
rect 483 1829 489 1834
rect 593 1828 599 1833
rect 703 1828 709 1833
rect 813 1828 819 1833
rect 1657 1889 1662 1897
rect 1653 1743 1661 1753
rect 920 1635 925 1643
rect 917 1617 925 1623
rect 1424 1657 1430 1663
rect 929 1446 935 1454
rect 1546 1463 1554 1480
rect 1658 1425 1662 1429
rect 1666 1425 1670 1429
rect 1674 1398 1682 1411
rect 53 1327 57 1333
rect 163 1326 167 1332
rect 273 1328 277 1334
rect 383 1326 387 1332
rect 493 1326 497 1332
rect 603 1326 607 1332
rect 713 1327 717 1333
rect 823 1326 827 1332
rect 904 1316 910 1320
rect 1424 1375 1430 1381
rect 1546 1316 1554 1333
rect 1654 1316 1658 1324
rect 1782 1264 1786 1268
rect 981 1218 991 1226
rect 1782 1189 1786 1193
rect 921 1181 925 1185
rect 12 1022 20 1039
rect 995 1161 1001 1167
rect 1105 1163 1111 1168
rect 1216 1164 1222 1168
rect 1327 1164 1333 1169
rect 1751 1135 1755 1139
rect 1750 1105 1754 1112
rect 1772 1097 1779 1101
rect 979 1044 987 1052
rect 979 1028 987 1036
rect 1744 1028 1752 1036
rect 1804 1264 1808 1268
rect 1789 1097 1793 1101
rect 1796 1256 1800 1260
rect 1762 1028 1770 1036
rect 1796 1024 1800 1028
rect 1804 1024 1808 1028
rect 1812 1158 1816 1162
rect 1812 1024 1816 1028
rect 1820 1024 1824 1028
rect 1828 1105 1836 1112
rect 1828 1024 1836 1028
rect 1844 1024 1852 1028
rect 156 1004 160 1010
rect 266 1003 270 1009
rect 376 1004 380 1010
rect 486 1003 490 1009
rect 596 1005 600 1011
rect 706 1004 710 1010
rect 816 1004 820 1010
rect 1796 745 1800 753
rect 1804 727 1808 733
rect 87 529 95 535
rect 189 529 197 535
rect 315 529 323 535
rect 417 529 425 535
rect 518 529 526 535
rect 645 529 653 535
rect 746 529 754 535
rect 848 529 856 535
rect 949 529 957 535
rect 1076 529 1084 535
rect 1177 529 1185 535
rect 1279 529 1287 535
rect 1405 529 1413 535
rect 1507 529 1515 535
rect 1622 529 1630 535
rect 1737 529 1745 535
rect 1812 493 1816 501
rect 1790 462 1794 466
rect 1820 462 1824 469
rect 45 428 51 434
rect 155 427 161 433
rect 265 425 271 431
rect 374 427 380 433
rect 485 427 491 433
rect 595 426 601 432
rect 705 427 711 433
rect 815 426 821 432
rect 925 426 931 432
rect 1035 428 1041 434
rect 1145 428 1151 434
rect 1255 427 1261 433
rect 1365 426 1371 432
rect 1475 427 1481 433
rect 1585 428 1591 434
rect 1695 426 1701 432
rect 1798 267 1806 277
rect 1817 123 1823 131
rect 1801 25 1807 31
rect 81 11 94 17
rect 191 11 204 17
rect 301 11 314 17
rect 411 11 424 17
rect 521 11 534 17
rect 631 11 644 17
rect 741 11 754 17
rect 851 11 864 17
rect 961 11 974 17
rect 1071 11 1084 17
rect 1181 11 1194 17
rect 1291 11 1304 17
rect 1401 11 1414 17
rect 1511 11 1524 17
rect 1621 11 1634 17
rect 1731 11 1744 17
<< psubstratepcontact >>
rect 1882 2006 1886 2014
rect 1950 2006 1954 2015
rect 1882 1981 1886 1989
rect 1950 1981 1954 1990
rect 1882 1956 1886 1964
rect 1950 1956 1954 1965
rect 1882 1931 1886 1939
rect 1950 1931 1954 1940
rect 1882 1906 1886 1914
rect 1950 1906 1954 1915
rect 1882 1881 1886 1889
rect 1950 1881 1954 1890
rect 1882 1856 1886 1864
rect 1950 1856 1954 1865
rect 1882 1831 1886 1839
rect 1950 1831 1954 1840
rect 1882 1806 1886 1814
rect 1950 1806 1954 1815
rect 1882 1781 1886 1789
rect 1950 1781 1954 1790
rect 1882 1756 1886 1764
rect 1950 1756 1954 1765
rect 1882 1731 1886 1739
rect 1950 1731 1954 1740
rect 1882 1706 1886 1714
rect 1950 1706 1954 1715
rect 1882 1681 1886 1689
rect 1950 1681 1954 1690
rect 1882 1656 1886 1664
rect 1950 1656 1954 1665
rect 1882 1631 1886 1639
rect 1950 1631 1954 1640
rect 1882 1606 1886 1614
rect 1950 1606 1954 1615
rect 1882 1581 1886 1589
rect 1950 1581 1954 1590
rect 1882 1556 1886 1564
rect 1950 1556 1954 1565
rect 1882 1531 1886 1539
rect 1950 1531 1954 1540
rect 1882 1506 1886 1514
rect 1950 1506 1954 1515
rect 1882 1481 1886 1489
rect 1950 1481 1954 1490
rect 1882 1456 1886 1464
rect 1950 1456 1954 1465
rect 1882 1431 1886 1439
rect 1950 1431 1954 1440
rect 1882 1406 1886 1414
rect 1950 1406 1954 1415
rect 1882 1381 1886 1389
rect 1950 1381 1954 1390
rect 1882 1356 1886 1364
rect 1950 1356 1954 1365
rect 1882 1331 1886 1339
rect 1950 1331 1954 1340
rect 1882 1306 1886 1314
rect 1950 1306 1954 1315
rect 1882 1281 1886 1289
rect 1950 1281 1954 1290
rect 1882 1256 1886 1264
rect 1950 1256 1954 1265
rect 1882 1231 1886 1239
rect 1950 1231 1954 1240
rect 1882 1206 1886 1214
rect 1950 1206 1954 1215
rect 1882 1181 1886 1189
rect 1950 1181 1954 1190
rect 1882 1156 1886 1164
rect 1950 1156 1954 1165
rect 1882 1131 1886 1139
rect 1950 1131 1954 1140
rect 1882 1106 1886 1114
rect 1950 1106 1954 1115
rect 1882 1081 1886 1089
rect 1950 1081 1954 1090
rect 1882 1056 1886 1064
rect 1950 1056 1954 1065
rect 1882 1031 1886 1039
rect 1950 1031 1954 1040
rect 1882 1006 1886 1014
rect 1950 1006 1954 1015
rect 1882 981 1886 989
rect 1950 981 1954 990
rect 1882 956 1886 964
rect 1950 956 1954 965
rect 1882 931 1886 939
rect 1950 931 1954 940
rect 1882 906 1886 914
rect 1950 906 1954 915
rect 1882 881 1886 889
rect 1950 881 1954 890
rect 1882 856 1886 864
rect 1950 856 1954 865
rect 1882 831 1886 839
rect 1950 831 1954 840
rect 1882 806 1886 814
rect 1950 806 1954 815
rect 1882 781 1886 789
rect 1950 781 1954 790
rect 1882 756 1886 764
rect 1950 756 1954 765
rect 1882 731 1886 739
rect 1950 731 1954 740
rect 1882 706 1886 714
rect 1950 706 1954 715
rect 1882 681 1886 689
rect 1950 681 1954 690
rect 1882 656 1886 664
rect 1950 656 1954 665
rect 1882 631 1886 639
rect 1950 631 1954 640
rect 1882 606 1886 614
rect 1950 606 1954 615
rect 1882 581 1886 589
rect 1950 581 1954 590
rect 1882 556 1886 564
rect 1950 556 1954 565
rect 1882 531 1886 539
rect 1950 531 1954 540
rect 1882 506 1886 514
rect 1950 506 1954 515
rect 1882 481 1886 489
rect 1950 481 1954 490
rect 1882 456 1886 464
rect 1950 456 1954 465
rect 1882 431 1886 439
rect 1950 431 1954 440
rect 1882 406 1886 414
rect 1950 406 1954 415
rect 1882 381 1886 389
rect 1950 381 1954 390
rect 1882 356 1886 364
rect 1950 356 1954 365
rect 1882 331 1886 339
rect 1950 331 1954 340
rect 1882 306 1886 314
rect 1950 306 1954 315
rect 1882 281 1886 289
rect 1950 281 1954 290
rect 1882 256 1886 264
rect 1950 256 1954 265
rect 1882 231 1886 239
rect 1950 231 1954 240
rect 1882 206 1886 214
rect 1950 206 1954 215
rect 1882 181 1886 189
rect 1950 181 1954 190
rect 1882 156 1886 164
rect 1950 156 1954 165
rect 1882 131 1886 139
rect 1950 131 1954 140
rect 1882 106 1886 114
rect 1950 106 1954 115
rect 1882 81 1886 89
rect 1950 81 1954 90
rect 1882 56 1886 64
rect 1950 56 1954 65
rect 1882 31 1886 39
rect 1950 31 1954 40
<< nsubstratencontact >>
rect 1916 2006 1920 2015
rect 1984 2006 1988 2015
rect 1916 1981 1920 1990
rect 1984 1981 1988 1990
rect 1916 1956 1920 1965
rect 1984 1956 1988 1965
rect 1916 1931 1920 1940
rect 1984 1931 1988 1940
rect 1916 1906 1920 1915
rect 1984 1906 1988 1915
rect 1916 1881 1920 1890
rect 1984 1881 1988 1890
rect 1916 1856 1920 1865
rect 1984 1856 1988 1865
rect 1916 1831 1920 1840
rect 1984 1831 1988 1840
rect 1916 1806 1920 1815
rect 1984 1806 1988 1815
rect 1916 1781 1920 1790
rect 1984 1781 1988 1790
rect 1916 1756 1920 1765
rect 1984 1756 1988 1765
rect 1916 1731 1920 1740
rect 1984 1731 1988 1740
rect 1916 1706 1920 1715
rect 1984 1706 1988 1715
rect 1916 1681 1920 1690
rect 1984 1681 1988 1690
rect 1916 1656 1920 1665
rect 1984 1656 1988 1665
rect 1916 1631 1920 1640
rect 1984 1631 1988 1640
rect 1916 1606 1920 1615
rect 1984 1606 1988 1615
rect 1916 1581 1920 1590
rect 1984 1581 1988 1590
rect 1916 1556 1920 1565
rect 1984 1556 1988 1565
rect 1916 1531 1920 1540
rect 1984 1531 1988 1540
rect 1916 1506 1920 1515
rect 1984 1506 1988 1515
rect 1916 1481 1920 1490
rect 1984 1481 1988 1490
rect 1916 1456 1920 1465
rect 1984 1456 1988 1465
rect 1916 1431 1920 1440
rect 1984 1431 1988 1440
rect 1916 1406 1920 1415
rect 1984 1406 1988 1415
rect 1916 1381 1920 1390
rect 1984 1381 1988 1390
rect 1916 1356 1920 1365
rect 1984 1356 1988 1365
rect 1916 1331 1920 1340
rect 1984 1331 1988 1340
rect 1916 1306 1920 1315
rect 1984 1306 1988 1315
rect 1916 1281 1920 1290
rect 1984 1281 1988 1290
rect 1916 1256 1920 1265
rect 1984 1256 1988 1265
rect 1916 1231 1920 1240
rect 1984 1231 1988 1240
rect 1916 1206 1920 1215
rect 1984 1206 1988 1215
rect 1916 1181 1920 1190
rect 1984 1181 1988 1190
rect 1916 1156 1920 1165
rect 1984 1156 1988 1165
rect 1916 1131 1920 1140
rect 1984 1131 1988 1140
rect 1916 1106 1920 1115
rect 1984 1106 1988 1115
rect 1916 1081 1920 1090
rect 1984 1081 1988 1090
rect 1916 1056 1920 1065
rect 1984 1056 1988 1065
rect 1916 1031 1920 1040
rect 1984 1031 1988 1040
rect 1916 1006 1920 1015
rect 1984 1006 1988 1015
rect 1916 981 1920 990
rect 1984 981 1988 990
rect 1916 956 1920 965
rect 1984 956 1988 965
rect 1916 931 1920 940
rect 1984 931 1988 940
rect 1916 906 1920 915
rect 1984 906 1988 915
rect 1916 881 1920 890
rect 1984 881 1988 890
rect 1916 856 1920 865
rect 1984 856 1988 865
rect 1916 831 1920 840
rect 1984 831 1988 840
rect 1916 806 1920 815
rect 1984 806 1988 815
rect 1916 781 1920 790
rect 1984 781 1988 790
rect 1916 756 1920 765
rect 1984 756 1988 765
rect 1916 731 1920 740
rect 1984 731 1988 740
rect 1916 706 1920 715
rect 1984 706 1988 715
rect 1916 681 1920 690
rect 1984 681 1988 690
rect 1916 656 1920 665
rect 1984 656 1988 665
rect 1916 631 1920 640
rect 1984 631 1988 640
rect 1916 606 1920 615
rect 1984 606 1988 615
rect 1916 581 1920 590
rect 1984 581 1988 590
rect 1916 556 1920 565
rect 1984 556 1988 565
rect 1916 531 1920 540
rect 1984 531 1988 540
rect 1916 506 1920 515
rect 1984 506 1988 515
rect 1916 481 1920 490
rect 1984 481 1988 490
rect 1916 456 1920 465
rect 1984 456 1988 465
rect 1916 431 1920 440
rect 1984 431 1988 440
rect 1916 406 1920 415
rect 1984 406 1988 415
rect 1916 381 1920 390
rect 1984 381 1988 390
rect 1916 356 1920 365
rect 1984 356 1988 365
rect 1916 331 1920 340
rect 1984 331 1988 340
rect 1916 306 1920 315
rect 1984 306 1988 315
rect 1916 281 1920 290
rect 1984 281 1988 290
rect 1916 256 1920 265
rect 1984 256 1988 265
rect 1916 231 1920 240
rect 1984 231 1988 240
rect 1916 206 1920 215
rect 1984 206 1988 215
rect 1916 181 1920 190
rect 1984 181 1988 190
rect 1916 156 1920 165
rect 1984 156 1988 165
rect 1916 131 1920 140
rect 1984 131 1988 140
rect 1916 106 1920 115
rect 1984 106 1988 115
rect 1916 81 1920 90
rect 1984 81 1988 90
rect 1916 56 1920 65
rect 1984 56 1988 65
rect 1916 31 1920 40
rect 1984 31 1988 40
use datapathL  datapathL_0
array 0 7 110 0 0 1803
timestamp 1428890255
transform 1 0 30 0 1 562
box 0 -542 110 1261
use rego  rego_2
timestamp 1428793378
transform 1 0 993 0 -1 1840
box 0 -160 110 279
use rego  rego_3
timestamp 1428793378
transform 1 0 1103 0 -1 1840
box 0 -160 110 279
use rego  rego_5
timestamp 1428793378
transform 1 0 1213 0 -1 1840
box 0 -160 110 279
use rego  rego_6
timestamp 1428793378
transform 1 0 1323 0 -1 1840
box 0 -160 110 279
use rego  rego_7
timestamp 1428793378
transform 1 0 1433 0 -1 1840
box 0 -160 110 279
use rego  rego_8
timestamp 1428793378
transform 1 0 1543 0 -1 1840
box 0 -160 110 279
use rego  rego_4
timestamp 1428793378
transform 1 0 993 0 1 1275
box 0 -160 110 279
use rego  rego_9
timestamp 1428793378
transform 1 0 1103 0 1 1275
box 0 -160 110 279
use rego  rego_1
timestamp 1428793378
transform 1 0 1213 0 1 1275
box 0 -160 110 279
use rego  rego_0
timestamp 1428793378
transform 1 0 1323 0 1 1275
box 0 -160 110 279
use and  and_0
timestamp 1427941063
transform 1 0 1736 0 1 1385
box -25 -23 14 33
use smlogic  smlogic_0
timestamp 1428811646
transform 1 0 1304 0 1 1193
box 123 -143 548 366
use datapathS  datapathS_0
array 0 7 110 0 0 974
timestamp 1428882048
transform 1 0 910 0 1 562
box 0 -542 110 432
<< labels >>
rlabel metal2 1790 495 1815 499 0 INBIT
rlabel metal1 -34 20 4 1822 0 Vdd
rlabel metal1 1828 19 1865 1021 0 GND
rlabel metal2 920 1643 928 2006 1 clk
rlabel space 1753 1119 1766 1121 1 start
rlabel metal2 1751 1135 1865 1139 1 start
rlabel metal1 1844 1028 1852 1344 1 reset
rlabel space 813 1785 819 1864 1 divisorin_0
rlabel m2contact 813 1828 819 1833 1 divisorin_0
rlabel m2contact 703 1828 709 1833 1 divisorin_1
rlabel m2contact 593 1828 599 1833 1 divisorin_2
rlabel m2contact 483 1829 489 1834 1 divisorin_3
rlabel m2contact 373 1829 379 1834 1 divisorin_4
rlabel m2contact 263 1828 269 1833 1 divisorin_5
rlabel m2contact 153 1829 159 1834 1 divisorin_6
rlabel metal2 1774 1032 1869 1036 1 dividendin_0
rlabel metal2 1665 1040 1869 1044 1 dividendin_1
rlabel metal2 1555 1048 1869 1052 1 dividendin_2
rlabel metal2 1445 1056 1869 1060 1 dividendin_3
rlabel metal2 1335 1064 1869 1068 1 dividendin_4
rlabel metal2 1225 1072 1869 1076 1 dividendin_5
rlabel metal2 1115 1080 1869 1084 1 dividendin_6
rlabel metal2 1005 1088 1869 1092 1 dividendin_7
rlabel space 1731 -21 1744 46 1 quotient_0
rlabel m2contact 1731 11 1744 17 1 quotient_0
rlabel m2contact 1621 11 1634 17 1 quotient_1
rlabel m2contact 1511 11 1524 17 1 quotient_2
rlabel m2contact 1401 11 1414 17 1 quotient_3
rlabel m2contact 1291 11 1304 17 1 quotient_4
rlabel m2contact 1181 11 1194 17 1 quotient_5
rlabel m2contact 1071 11 1084 17 1 quotient_6
rlabel m2contact 961 11 974 17 1 quotient_7
rlabel m2contact 81 11 94 17 1 remainder_6
rlabel m2contact 191 11 204 17 1 remainder_5
rlabel m2contact 301 11 314 17 1 remainder_4
rlabel m2contact 411 11 424 17 1 remainder_3
rlabel m2contact 521 11 534 17 1 remainder_2
rlabel m2contact 631 11 644 17 1 remainder_1
rlabel m2contact 741 11 754 17 1 remainder_0
rlabel space 1740 1329 1742 1370 1 SB1
rlabel polysilicon 1740 1410 1742 1434 1 SB1
rlabel polysilicon 1730 1410 1732 1434 1 SB0
rlabel polysilicon 1707 1433 1715 1434 1 sign
rlabel space 1613 1113 1651 1115 1 SB0_out
rlabel metal2 917 1328 925 1617 1 clkload
rlabel space 1666 1342 1670 1559 1 nextsb1
rlabel m2contact 1666 1425 1670 1429 1 nextsb1
rlabel m2contact 1658 1425 1662 1429 1 nextsb0
rlabel m2contact 816 1004 820 1010 1 sum0
rlabel m2contact 706 1004 710 1010 1 sum1
rlabel m2contact 596 1005 600 1011 1 sum2
rlabel m2contact 486 1003 490 1009 1 sum3
rlabel m2contact 376 1004 380 1010 1 sum4
rlabel space 266 989 270 1021 1 sum5
rlabel space 156 989 160 1021 1 sum6
rlabel m2contact 266 1003 270 1009 1 sum5
rlabel m2contact 156 1004 160 1010 1 sum6
rlabel m2contact 823 1326 827 1332 1 divregout0
rlabel m2contact 713 1327 717 1333 1 divregout1
rlabel m2contact 603 1326 607 1332 1 divregout2
rlabel m2contact 493 1326 497 1332 1 divregout3
rlabel m2contact 383 1326 387 1332 1 divregout4
rlabel m2contact 273 1328 277 1334 1 divregout5
rlabel m2contact 163 1326 167 1332 1 divregout6
rlabel m2contact 53 1327 57 1333 1 divregout7
rlabel m2contact 1737 529 1745 535 1 qmuxout0
rlabel m2contact 1622 529 1630 535 1 qmuxout1
rlabel m2contact 1507 529 1515 535 1 qmuxout2
rlabel m2contact 1405 529 1413 535 1 qmuxout3
rlabel m2contact 1279 529 1287 535 1 qmuxout4
rlabel m2contact 1177 529 1185 535 1 qmuxout5
rlabel m2contact 1076 529 1084 535 1 qmuxout6
rlabel m2contact 949 529 957 535 1 qmuxout7
rlabel m2contact 746 529 754 535 1 rmuxout1
rlabel m2contact 645 529 653 535 1 rmuxout2
rlabel m2contact 518 529 526 535 1 rmuxout3
rlabel m2contact 417 529 425 535 1 rmuxout4
rlabel m2contact 315 529 323 535 1 rmuxout5
rlabel m2contact 189 529 197 535 1 rmuxout6
rlabel m2contact 87 529 95 535 1 rmuxout7
rlabel metal1 1775 1314 1812 1318 1 shift
rlabel metal1 1775 1291 1789 1295 1 load
rlabel metal2 1786 1264 1804 1268 1 sel1
rlabel metal1 1796 1024 1800 1252 1 sel0
rlabel space 1776 1189 1782 1193 1 add
rlabel metal2 1778 1158 1812 1162 1 inbit
rlabel m2contact 1782 1189 1786 1193 1 add
rlabel m2contact 1327 1164 1333 1169 1 validregs0
rlabel m2contact 1216 1164 1222 1168 1 validregs1
rlabel m2contact 1105 1163 1111 1168 1 validregs2
rlabel m2contact 995 1161 1001 1167 1 validregs3
rlabel space 1011 1952 1024 1957 1 validregs4
rlabel metal2 1104 1599 1110 2017 1 validregs4
rlabel metal2 1214 1599 1220 2017 1 validregs5
rlabel metal2 1324 1599 1330 2017 1 validregs6
rlabel metal2 1434 1599 1440 2017 1 validregs7
rlabel space 1695 421 1701 457 1 qregin
rlabel m2contact 925 426 931 432 1 qregin7
rlabel m2contact 1035 428 1041 434 1 qregin6
rlabel m2contact 1145 428 1151 434 1 qregin5
rlabel m2contact 1255 427 1261 433 1 qregin4
rlabel m2contact 1365 426 1371 432 1 qregin3
rlabel m2contact 1475 427 1481 433 1 qregin2
rlabel m2contact 1585 428 1591 434 1 qregin1
rlabel m2contact 45 428 51 434 1 rregin7
rlabel m2contact 155 427 161 433 1 rregin6
rlabel m2contact 265 425 271 431 1 rregin5
rlabel m2contact 374 427 380 433 1 rregin4
rlabel m2contact 485 427 491 433 1 rregin3
rlabel m2contact 595 426 601 432 1 rregin2
rlabel m2contact 705 427 711 433 1 rregin1
rlabel m2contact 815 426 821 432 1 rregin0
rlabel metal2 1451 2012 1550 2017 1 valid
rlabel m2contact 1695 426 1701 432 1 qregin0
rlabel m2contact 848 529 856 535 1 rmuxout0
<< end >>
