magic
tech scmos
timestamp 1428801662
<< pwell >>
rect 0 240 110 279
rect 0 95 110 151
rect 0 -109 110 -24
<< nwell >>
rect 0 157 110 234
rect 0 -18 110 89
rect 0 -160 110 -113
<< polysilicon >>
rect 22 250 24 252
rect 34 250 60 252
rect 56 248 60 250
rect 74 250 77 252
rect 87 250 101 252
rect 56 225 64 248
rect 22 223 24 225
rect 44 223 53 225
rect 56 223 67 225
rect 87 223 89 225
rect 48 214 53 223
rect 48 208 58 214
rect 22 184 24 186
rect 74 184 76 186
rect 22 162 24 164
rect 74 162 76 164
rect 11 160 24 162
rect 18 150 24 160
rect 11 148 24 150
rect 54 160 76 162
rect 61 150 76 160
rect 54 148 76 150
rect 22 146 24 148
rect 74 146 76 148
rect 22 134 24 136
rect 74 134 76 136
rect 45 111 47 113
rect 82 111 84 113
rect 45 99 47 101
rect 45 97 62 99
rect 45 87 55 97
rect 45 85 62 87
rect 82 97 84 101
rect 82 95 107 97
rect 82 89 94 95
rect 82 87 107 89
rect 45 83 47 85
rect 82 83 84 87
rect 45 61 47 63
rect 82 61 84 63
rect 64 39 87 43
rect 64 37 66 39
rect 72 37 74 39
rect 15 30 22 36
rect 15 1 19 30
rect 21 17 23 19
rect 43 17 52 19
rect 82 33 87 39
rect 94 37 96 39
rect 15 -1 23 1
rect 43 -1 45 1
rect 15 -40 22 -1
rect 48 -18 52 17
rect 64 16 66 18
rect 72 16 74 18
rect 64 7 66 9
rect 72 7 74 9
rect 64 -15 66 -13
rect 72 -15 74 -13
rect 82 -15 87 22
rect 94 15 96 17
rect 94 12 109 15
rect 94 8 96 10
rect 64 -16 87 -15
rect 94 -16 96 -12
rect 64 -18 96 -16
rect 37 -21 52 -18
rect 48 -22 52 -21
rect 49 -30 52 -22
rect 25 -32 27 -30
rect 37 -32 52 -30
rect 82 -26 96 -18
rect 15 -42 25 -40
rect 23 -48 25 -42
rect 63 -45 65 -43
rect 71 -45 73 -43
rect 23 -50 27 -48
rect 37 -50 39 -48
rect 82 -49 87 -26
rect 94 -28 96 -26
rect 94 -40 96 -38
rect 104 -42 109 12
rect 94 -46 109 -42
rect 94 -48 96 -46
rect 104 -49 109 -46
rect 63 -66 65 -65
rect 71 -66 73 -65
rect 94 -66 96 -58
rect 63 -68 96 -66
rect 65 -90 67 -88
rect 93 -90 95 -88
rect 8 -99 10 -97
rect 40 -99 48 -97
rect 43 -117 48 -99
rect 65 -102 67 -100
rect 93 -102 95 -100
rect 65 -104 79 -102
rect 93 -104 106 -102
rect 65 -114 72 -104
rect 97 -106 106 -104
rect 97 -112 99 -106
rect 97 -114 106 -112
rect 65 -116 79 -114
rect 93 -116 106 -114
rect 43 -126 52 -117
rect 8 -128 10 -126
rect 40 -127 52 -126
rect 65 -118 67 -116
rect 93 -118 95 -116
rect 40 -128 48 -127
rect 43 -134 48 -128
rect 8 -136 10 -134
rect 40 -136 48 -134
rect 65 -140 67 -138
rect 93 -140 95 -138
<< ndiffusion >>
rect 24 252 34 253
rect 24 249 34 250
rect 77 252 87 253
rect 77 249 87 250
rect 21 136 22 146
rect 24 136 25 146
rect 73 136 74 146
rect 76 136 77 146
rect 44 101 45 111
rect 47 101 48 111
rect 81 101 82 111
rect 84 101 85 111
rect 27 -30 37 -29
rect 27 -33 37 -32
rect 27 -48 37 -47
rect 27 -51 37 -50
rect 58 -65 63 -45
rect 65 -65 71 -45
rect 73 -65 78 -45
rect 93 -38 94 -28
rect 96 -38 97 -28
rect 93 -58 94 -48
rect 96 -58 97 -48
rect 10 -97 40 -96
rect 10 -100 40 -99
rect 64 -100 65 -90
rect 67 -100 68 -90
rect 92 -100 93 -90
rect 95 -100 96 -90
<< pdiffusion >>
rect 24 225 44 226
rect 67 225 87 226
rect 24 222 44 223
rect 67 222 87 223
rect 21 164 22 184
rect 24 164 25 184
rect 73 164 74 184
rect 76 164 77 184
rect 44 63 45 83
rect 47 63 48 83
rect 81 63 82 83
rect 84 63 85 83
rect 23 19 43 20
rect 63 18 64 37
rect 66 18 67 37
rect 71 18 72 37
rect 74 18 75 37
rect 23 16 43 17
rect 23 1 43 2
rect 23 -2 43 -1
rect 63 -13 64 7
rect 66 -13 67 7
rect 71 -13 72 7
rect 74 -13 75 7
rect 93 17 94 37
rect 96 17 97 37
rect 93 -12 94 8
rect 96 -12 97 8
rect 10 -126 40 -125
rect 10 -129 40 -128
rect 10 -134 40 -133
rect 10 -137 40 -136
rect 64 -138 65 -118
rect 67 -138 68 -118
rect 92 -138 93 -118
rect 95 -138 96 -118
<< metal1 >>
rect 0 277 110 279
rect 0 265 14 277
rect 21 265 42 277
rect 49 265 71 277
rect 78 265 110 277
rect 0 263 110 265
rect 13 253 24 257
rect 13 241 21 253
rect 13 235 15 241
rect 13 222 21 235
rect 49 248 60 254
rect 87 253 97 257
rect 24 241 87 245
rect 24 235 28 241
rect 34 235 87 241
rect 24 230 87 235
rect 90 240 97 253
rect 96 234 97 240
rect 90 222 97 234
rect 13 218 24 222
rect 87 218 97 222
rect 64 209 69 214
rect 101 214 107 248
rect 75 209 107 214
rect 64 208 107 209
rect 0 203 110 205
rect 0 191 16 203
rect 23 191 41 203
rect 48 191 79 203
rect 86 191 110 203
rect 0 189 110 191
rect 13 184 21 189
rect 65 184 73 189
rect 13 164 17 184
rect 29 164 49 184
rect 65 164 69 184
rect 81 164 98 184
rect 37 162 49 164
rect 37 160 61 162
rect 18 158 33 160
rect 18 152 27 158
rect 18 150 33 152
rect 37 150 54 160
rect 37 148 61 150
rect 86 159 98 164
rect 86 153 87 159
rect 93 153 98 159
rect 37 146 49 148
rect 86 146 98 153
rect 13 136 17 146
rect 29 145 49 146
rect 29 138 33 145
rect 40 138 49 145
rect 29 136 49 138
rect 65 136 69 146
rect 81 136 98 146
rect 13 131 21 136
rect 65 131 73 136
rect 0 129 110 131
rect 0 117 14 129
rect 21 117 42 129
rect 49 117 71 129
rect 78 117 110 129
rect 0 115 110 117
rect 48 111 56 115
rect 85 111 93 115
rect 35 97 40 111
rect 52 101 56 111
rect 62 101 77 111
rect 89 101 93 111
rect 0 95 40 97
rect 0 88 36 95
rect 0 87 40 88
rect 25 63 40 87
rect 62 83 74 101
rect 100 95 110 97
rect 107 89 110 95
rect 100 87 110 89
rect 52 63 56 83
rect 62 74 77 83
rect 67 67 77 74
rect 62 63 77 67
rect 89 63 93 83
rect 48 57 56 63
rect 85 57 93 63
rect 0 55 110 57
rect 0 44 16 55
rect 23 44 41 55
rect 48 44 79 55
rect 86 44 110 55
rect 0 41 110 44
rect 67 37 71 41
rect 97 37 101 41
rect 30 30 35 36
rect 10 24 59 27
rect 10 20 23 24
rect 43 20 59 24
rect 10 -36 16 20
rect 56 18 59 20
rect 56 15 63 18
rect 23 7 54 12
rect 67 7 71 18
rect 75 15 79 18
rect 82 33 89 37
rect 87 22 89 33
rect 82 17 89 22
rect 97 8 101 17
rect 23 6 59 7
rect 43 2 59 6
rect 22 -6 23 -2
rect 22 -13 27 -6
rect 46 -9 50 2
rect 22 -20 23 -13
rect 22 -29 27 -20
rect 31 -16 37 -15
rect 40 -13 50 -9
rect 10 -41 22 -36
rect 0 -57 11 -49
rect 14 -51 22 -41
rect 40 -37 44 -13
rect 59 -16 63 -13
rect 75 -16 79 -13
rect 59 -20 79 -16
rect 84 -23 89 8
rect 47 -27 89 -23
rect 27 -43 40 -37
rect 14 -55 27 -51
rect 37 -55 41 -51
rect 5 -59 11 -57
rect 48 -59 52 -27
rect 5 -67 52 -59
rect 58 -34 67 -30
rect 71 -34 78 -30
rect 84 -34 89 -27
rect 58 -65 62 -34
rect 66 -70 70 -45
rect 74 -65 78 -34
rect 97 -48 101 -38
rect 82 -49 89 -48
rect 87 -57 89 -49
rect 82 -58 89 -57
rect 97 -70 101 -58
rect 0 -72 110 -70
rect 0 -84 14 -72
rect 21 -84 42 -72
rect 49 -84 71 -72
rect 78 -84 110 -72
rect 0 -86 110 -84
rect 10 -92 40 -86
rect 68 -90 76 -86
rect 96 -90 104 -86
rect 2 -104 10 -100
rect 2 -112 40 -104
rect 2 -114 18 -112
rect 2 -129 7 -114
rect 31 -114 40 -112
rect 55 -107 60 -90
rect 72 -100 76 -90
rect 79 -100 88 -90
rect 100 -100 104 -90
rect 55 -117 60 -113
rect 40 -125 48 -121
rect 2 -133 10 -129
rect 43 -137 48 -125
rect 56 -127 60 -117
rect 79 -118 83 -100
rect 94 -112 99 -106
rect 40 -141 48 -137
rect 55 -138 60 -127
rect 72 -138 76 -118
rect 79 -132 88 -118
rect 85 -138 88 -132
rect 100 -138 104 -118
rect 10 -144 48 -141
rect 68 -144 76 -138
rect 96 -144 104 -138
rect 0 -146 110 -144
rect 0 -158 16 -146
rect 23 -158 41 -146
rect 48 -158 79 -146
rect 86 -158 110 -146
rect 0 -160 110 -158
<< metal2 >>
rect 15 241 21 277
rect 46 260 56 261
rect 46 254 49 260
rect 55 254 56 260
rect 25 241 36 242
rect 25 235 28 241
rect 34 235 36 241
rect 25 158 36 235
rect 25 152 27 158
rect 33 152 36 158
rect 25 151 36 152
rect 14 145 40 147
rect 14 138 33 145
rect 14 136 40 138
rect 14 -11 21 136
rect 46 122 56 254
rect 85 234 90 240
rect 25 115 56 122
rect 64 209 69 215
rect 25 74 32 115
rect 64 108 75 209
rect 85 159 96 234
rect 85 153 87 159
rect 93 153 103 159
rect 85 151 103 153
rect 64 103 79 108
rect 71 95 79 103
rect 43 88 79 95
rect 25 67 60 74
rect 25 36 32 67
rect 71 54 79 88
rect 46 47 79 54
rect 25 30 35 36
rect 25 29 41 30
rect 46 25 52 47
rect 31 21 52 25
rect 31 -9 37 21
rect 75 1 79 10
rect 14 -13 27 -11
rect 14 -20 23 -13
rect 54 -4 79 1
rect 54 -19 58 -4
rect 27 -20 58 -19
rect 14 -22 58 -20
rect 23 -23 58 -22
rect 99 -23 103 151
rect 67 -27 106 -23
rect 67 -30 71 -27
rect 44 -38 63 -37
rect 44 -43 74 -38
rect 45 -55 61 -51
rect 51 -107 61 -55
rect 66 -65 74 -43
rect 66 -73 95 -65
rect 51 -113 55 -107
rect 87 -106 95 -73
rect 87 -112 88 -106
rect 94 -112 95 -106
rect 79 -132 88 -130
rect 85 -138 88 -132
rect 79 -148 88 -138
rect 51 -156 88 -148
rect 51 -160 64 -156
<< ntransistor >>
rect 24 250 34 252
rect 77 250 87 252
rect 22 136 24 146
rect 74 136 76 146
rect 45 101 47 111
rect 82 101 84 111
rect 27 -32 37 -30
rect 27 -50 37 -48
rect 63 -65 65 -45
rect 71 -65 73 -45
rect 94 -38 96 -28
rect 94 -58 96 -48
rect 10 -99 40 -97
rect 65 -100 67 -90
rect 93 -100 95 -90
<< ptransistor >>
rect 24 223 44 225
rect 67 223 87 225
rect 22 164 24 184
rect 74 164 76 184
rect 45 63 47 83
rect 82 63 84 83
rect 23 17 43 19
rect 64 18 66 37
rect 72 18 74 37
rect 23 -1 43 1
rect 64 -13 66 7
rect 72 -13 74 7
rect 94 17 96 37
rect 94 -12 96 8
rect 10 -128 40 -126
rect 10 -136 40 -134
rect 65 -138 67 -118
rect 93 -138 95 -118
<< polycontact >>
rect 60 248 66 254
rect 101 248 107 254
rect 58 208 64 214
rect 11 150 18 160
rect 54 150 61 160
rect 55 87 62 97
rect 94 89 107 95
rect 22 30 30 36
rect 82 22 87 33
rect 31 -22 37 -16
rect 82 -57 87 -49
rect 104 -57 110 -49
rect 72 -114 79 -104
rect 99 -112 106 -106
rect 52 -127 56 -117
<< ndcontact >>
rect 24 253 34 257
rect 24 245 34 249
rect 77 253 87 257
rect 77 245 87 249
rect 17 136 21 146
rect 25 136 29 146
rect 69 136 73 146
rect 77 136 81 146
rect 40 101 44 111
rect 48 101 52 111
rect 77 101 81 111
rect 85 101 89 111
rect 27 -29 37 -25
rect 27 -37 37 -33
rect 27 -47 37 -43
rect 27 -55 37 -51
rect 89 -38 93 -28
rect 97 -38 101 -28
rect 89 -58 93 -48
rect 97 -58 101 -48
rect 10 -96 40 -92
rect 10 -104 40 -100
rect 60 -100 64 -90
rect 68 -100 72 -90
rect 88 -100 92 -90
rect 96 -100 100 -90
<< pdcontact >>
rect 24 226 44 230
rect 67 226 87 230
rect 24 218 44 222
rect 67 218 87 222
rect 17 164 21 184
rect 25 164 29 184
rect 69 164 73 184
rect 77 164 81 184
rect 40 63 44 83
rect 48 63 52 83
rect 77 63 81 83
rect 85 63 89 83
rect 23 20 43 24
rect 59 18 63 37
rect 67 18 71 37
rect 75 18 79 37
rect 23 12 43 16
rect 23 2 43 6
rect 23 -6 43 -2
rect 59 -13 63 7
rect 67 -13 71 7
rect 75 -13 79 7
rect 89 17 93 37
rect 97 17 101 37
rect 89 -12 93 8
rect 97 -12 101 8
rect 10 -125 40 -121
rect 10 -133 40 -129
rect 10 -141 40 -137
rect 60 -138 64 -118
rect 68 -138 72 -118
rect 88 -138 92 -118
rect 96 -138 100 -118
<< m2contact >>
rect 49 254 55 260
rect 15 235 21 241
rect 28 235 34 241
rect 90 234 96 240
rect 69 209 75 215
rect 27 152 33 158
rect 87 153 93 159
rect 33 138 40 145
rect 36 88 43 95
rect 60 67 67 74
rect 35 30 41 36
rect 59 10 63 15
rect 75 10 79 15
rect 23 -20 27 -13
rect 31 -15 37 -9
rect 40 -43 44 -37
rect 41 -55 45 -51
rect 67 -34 71 -30
rect 18 -117 31 -112
rect 55 -113 61 -107
rect 88 -112 94 -106
rect 79 -138 85 -132
<< psubstratepcontact >>
rect 14 265 21 277
rect 42 265 49 277
rect 71 265 78 277
rect 14 117 21 129
rect 42 117 49 129
rect 71 117 78 129
rect 14 -84 21 -72
rect 42 -84 49 -72
rect 71 -84 78 -72
<< nsubstratencontact >>
rect 16 191 23 203
rect 41 191 48 203
rect 79 191 86 203
rect 16 44 23 55
rect 41 44 48 55
rect 79 44 86 55
rect 16 -158 23 -146
rect 41 -158 48 -146
rect 79 -158 86 -146
<< labels >>
rlabel metal1 37 148 54 162 0 REGMEM
rlabel metal1 62 74 74 111 0 INCLKn
rlabel metal1 25 63 40 97 0 INCLK
rlabel polysilicon 82 87 94 97 0 CLK
rlabel metal1 79 -138 88 -118 0 REGOUT
rlabel metal1 2 -114 18 -108 0 REGBUF
rlabel space 12 233 21 279 0 REGIN
rlabel polysilicon 104 -46 109 -26 0 RST
rlabel metal2 66 -73 74 -38 1 REGOUTn
rlabel space 592 -854 598 -818 8 qregin
<< end >>
