magic
tech scmos
timestamp 1428788720
<< pwell >>
rect 0 690 38 700
rect 6 684 38 690
rect 17 676 38 684
<< polysilicon >>
rect 0 185 4 189
<< metal1 >>
rect 1 1256 4 1257
rect 0 1249 4 1256
rect 1 1247 4 1249
rect 105 1176 110 1183
rect 0 1100 7 1107
rect 106 987 110 994
rect 0 859 7 866
rect 101 783 110 790
rect 0 659 8 666
rect 0 619 3 623
rect 103 555 110 562
rect 0 427 8 434
rect 103 322 110 329
rect 0 213 8 222
rect 0 166 3 170
rect 101 93 110 102
rect 0 -14 5 -5
rect 104 -50 110 -41
rect 0 -116 9 -107
rect 105 -189 110 -180
rect 0 -264 4 -255
rect 104 -338 110 -329
rect 0 -465 6 -456
rect 102 -540 110 -531
<< metal2 >>
rect 13 1254 19 1261
rect 27 781 54 788
rect 0 189 6 670
rect 16 427 65 432
rect 2 185 6 189
rect 0 -15 6 185
rect 0 -21 65 -15
rect 4 -493 10 -21
rect 96 -27 105 -15
rect 27 -33 105 -27
rect 27 -45 31 -33
rect 37 -105 41 -103
rect 21 -110 41 -105
rect 4 -500 31 -493
<< m2contact >>
rect 95 426 101 432
use reg  reg_0 ../cells
timestamp 1428788720
transform 1 0 18 0 1 982
box -18 -201 92 279
use adder  adder_0 ../cells
timestamp 1428734989
transform 1 0 0 0 1 432
box 0 0 110 356
use mux  mux_0 ../cells
timestamp 1428736483
transform 1 0 20 0 1 -15
box -20 0 90 447
use shifter  shifter_0 ../cells
timestamp 1428356401
transform 1 0 35 0 1 -106
box -35 3 75 68
use rego  rego_0 ../cells
timestamp 1428788278
transform 1 0 0 0 1 -382
box 0 -160 110 279
<< end >>
