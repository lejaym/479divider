magic
tech scmos
timestamp 1428354897
<< pwell >>
rect -18 242 92 279
rect -18 81 92 150
rect -18 -150 92 -66
<< nwell >>
rect -18 160 92 232
rect -18 -56 92 71
rect -18 -201 92 -150
<< polysilicon >>
rect -1 250 1 252
rect 11 250 14 252
rect 51 250 54 252
rect 64 250 83 252
rect -1 223 1 225
rect 21 223 27 225
rect 23 210 27 223
rect 75 225 83 250
rect 38 223 44 225
rect 64 223 66 225
rect 75 219 76 225
rect 82 219 83 225
rect 23 209 41 210
rect 23 206 49 209
rect 4 184 6 186
rect 56 184 58 186
rect 4 162 6 164
rect 56 162 58 164
rect -7 160 6 162
rect 0 150 6 160
rect -7 148 6 150
rect 36 160 58 162
rect 43 150 58 160
rect 36 148 58 150
rect 4 146 6 148
rect 56 146 58 148
rect 4 134 6 136
rect 56 134 58 136
rect 26 111 28 113
rect 64 111 66 113
rect 26 99 28 101
rect 64 99 66 101
rect -13 91 15 99
rect 26 95 51 99
rect 64 95 92 99
rect 26 91 28 93
rect 8 71 15 91
rect 26 79 28 81
rect 46 80 51 95
rect 64 91 66 93
rect 82 91 92 95
rect 26 78 40 79
rect 26 72 28 78
rect 26 71 40 72
rect 26 69 28 71
rect 49 70 51 80
rect 26 47 28 49
rect 46 45 51 70
rect 64 79 66 81
rect 64 73 74 79
rect 64 69 66 73
rect 64 47 66 49
rect 82 45 87 91
rect 26 42 51 45
rect 64 42 87 45
rect 26 40 28 42
rect 64 40 66 42
rect 26 18 28 20
rect 64 18 66 20
rect 47 -4 49 -2
rect 72 -4 74 -2
rect -3 -40 4 -5
rect 7 -24 9 -22
rect 29 -24 38 -22
rect -3 -42 9 -40
rect 29 -42 31 -40
rect -3 -81 4 -42
rect 33 -63 38 -24
rect 47 -45 49 -43
rect 58 -45 63 -19
rect 72 -26 74 -24
rect 72 -29 87 -26
rect 72 -33 74 -31
rect 47 -52 63 -45
rect 32 -71 38 -63
rect 7 -73 9 -71
rect 19 -73 38 -71
rect 58 -57 63 -52
rect 72 -57 74 -53
rect 58 -67 74 -57
rect -3 -83 7 -81
rect 5 -89 7 -83
rect 5 -91 9 -89
rect 19 -91 22 -89
rect 58 -90 63 -67
rect 72 -69 74 -67
rect 72 -81 74 -79
rect 82 -83 87 -29
rect 72 -87 87 -83
rect 72 -89 74 -87
rect 82 -90 87 -87
rect 72 -101 74 -99
rect 15 -131 17 -129
rect 57 -131 59 -129
rect 15 -143 17 -141
rect 57 -143 59 -141
rect 15 -145 32 -143
rect 15 -155 25 -145
rect 15 -157 32 -155
rect 57 -145 70 -143
rect 57 -155 63 -145
rect 57 -157 70 -155
rect 15 -159 17 -157
rect 57 -159 59 -157
rect 15 -181 17 -179
rect 57 -181 59 -179
<< ndiffusion >>
rect 1 252 11 253
rect 1 249 11 250
rect 54 252 64 253
rect 54 249 64 250
rect 3 136 4 146
rect 6 136 7 146
rect 55 136 56 146
rect 58 136 59 146
rect 25 101 26 111
rect 28 101 29 111
rect 63 101 64 111
rect 66 101 67 111
rect 25 81 26 91
rect 28 81 29 91
rect 63 81 64 91
rect 66 81 67 91
rect 9 -71 19 -70
rect 9 -74 19 -73
rect 9 -89 19 -88
rect 71 -79 72 -69
rect 74 -79 75 -69
rect 9 -92 19 -91
rect 71 -99 72 -89
rect 74 -99 75 -89
rect 14 -141 15 -131
rect 17 -141 18 -131
rect 56 -141 57 -131
rect 59 -141 60 -131
<< pdiffusion >>
rect 1 225 21 226
rect 1 222 21 223
rect 44 225 64 226
rect 44 222 64 223
rect 3 164 4 184
rect 6 164 7 184
rect 55 164 56 184
rect 58 164 59 184
rect 25 49 26 69
rect 28 49 29 69
rect 63 49 64 69
rect 66 49 67 69
rect 25 20 26 40
rect 28 20 29 40
rect 63 20 64 40
rect 66 20 67 40
rect 9 -22 29 -21
rect 9 -25 29 -24
rect 9 -40 29 -39
rect 9 -43 29 -42
rect 46 -43 47 -4
rect 49 -43 50 -4
rect 71 -24 72 -4
rect 74 -24 75 -4
rect 71 -53 72 -33
rect 74 -53 75 -33
rect 14 -179 15 -159
rect 17 -179 18 -159
rect 56 -179 57 -159
rect 59 -179 60 -159
<< metal1 >>
rect -18 277 92 279
rect -18 265 -4 277
rect 3 265 24 277
rect 31 265 53 277
rect 60 265 92 277
rect -18 263 92 265
rect -13 253 1 257
rect 14 256 30 257
rect 14 255 23 256
rect -13 241 -2 253
rect 20 250 23 255
rect 29 250 30 256
rect 64 253 77 257
rect 20 249 30 250
rect 5 241 64 245
rect -13 235 -5 241
rect 11 235 64 241
rect -13 222 -2 235
rect 5 230 64 235
rect -13 218 1 222
rect 29 221 32 227
rect 67 240 77 253
rect 73 234 77 240
rect 67 229 77 234
rect 67 222 73 229
rect 29 219 38 221
rect 35 213 38 219
rect 64 218 73 222
rect 82 219 83 225
rect 29 212 38 213
rect 47 209 50 215
rect 76 209 83 219
rect 41 208 56 209
rect -18 203 92 205
rect -18 191 -2 203
rect 5 191 23 203
rect 30 191 61 203
rect 68 191 92 203
rect -18 189 92 191
rect -5 184 3 189
rect 47 184 55 189
rect -5 164 -1 184
rect 11 164 31 184
rect 47 164 51 184
rect 19 162 31 164
rect 19 160 43 162
rect 0 157 15 160
rect 0 151 9 157
rect 0 150 15 151
rect 19 150 36 160
rect 63 159 72 184
rect 66 153 72 159
rect 19 148 43 150
rect 19 146 31 148
rect -5 136 -1 146
rect 11 145 31 146
rect 11 138 15 145
rect 22 138 31 145
rect 11 136 31 138
rect 47 136 51 146
rect 63 136 72 153
rect -5 131 3 136
rect 47 131 55 136
rect -18 129 92 131
rect -18 117 -4 129
rect 3 117 24 129
rect 31 117 53 129
rect 60 117 92 129
rect -18 115 92 117
rect 29 111 33 115
rect 67 111 71 115
rect -3 109 21 111
rect -3 103 12 109
rect 18 103 21 109
rect -3 101 21 103
rect -3 79 7 101
rect 29 91 33 101
rect -13 73 7 79
rect -3 40 7 73
rect 11 79 21 91
rect 36 101 59 111
rect 11 71 15 79
rect 36 78 42 101
rect 67 91 71 101
rect 40 72 42 78
rect 11 58 21 71
rect 17 52 21 58
rect 11 49 21 52
rect 29 40 33 49
rect -3 20 21 40
rect 36 40 42 72
rect 45 80 63 81
rect 49 77 63 80
rect 49 71 54 77
rect 60 71 63 77
rect 79 73 92 79
rect 49 70 63 71
rect 45 69 63 70
rect 67 40 71 49
rect 36 32 59 40
rect 36 26 39 32
rect 45 26 59 32
rect 36 20 59 26
rect 29 16 33 20
rect 67 16 71 20
rect -18 14 92 16
rect -18 3 -2 14
rect 5 3 23 14
rect 30 3 61 14
rect 68 3 92 14
rect -18 0 92 3
rect 50 -4 54 0
rect 75 -4 79 0
rect 12 -11 16 -5
rect -8 -21 9 -17
rect -8 -77 -2 -21
rect 29 -29 42 -25
rect 9 -35 42 -29
rect 29 -39 42 -35
rect 4 -47 9 -43
rect 4 -54 19 -47
rect 4 -61 10 -54
rect 17 -61 19 -54
rect 4 -66 19 -61
rect 4 -70 9 -66
rect 30 -57 32 -51
rect 24 -63 32 -57
rect 24 -71 27 -63
rect 35 -56 42 -39
rect 58 -8 67 -4
rect 63 -19 67 -8
rect 58 -24 67 -19
rect 75 -33 79 -24
rect 35 -63 54 -56
rect 35 -69 48 -63
rect -8 -82 4 -77
rect -4 -90 4 -82
rect 35 -78 42 -69
rect 62 -75 67 -33
rect 9 -84 42 -78
rect 46 -84 67 -75
rect -18 -98 -7 -90
rect 2 -92 4 -90
rect 2 -96 9 -92
rect -13 -100 -7 -98
rect 46 -100 54 -84
rect 75 -89 79 -79
rect 58 -90 67 -89
rect 63 -98 67 -90
rect 58 -99 67 -98
rect 88 -98 92 -90
rect -13 -108 54 -100
rect 75 -111 79 -99
rect -18 -113 92 -111
rect -18 -125 -4 -113
rect 3 -125 24 -113
rect 31 -125 53 -113
rect 60 -125 92 -113
rect -18 -127 92 -125
rect 18 -131 26 -127
rect 60 -131 68 -127
rect -7 -141 10 -131
rect 22 -141 26 -131
rect 32 -141 52 -131
rect 64 -141 68 -131
rect -7 -148 5 -141
rect -7 -154 -2 -148
rect 4 -154 5 -148
rect -7 -159 5 -154
rect 32 -159 44 -141
rect 48 -147 63 -145
rect 54 -153 63 -147
rect 48 -155 63 -153
rect -7 -179 10 -159
rect 22 -179 26 -159
rect 32 -168 52 -159
rect 32 -175 36 -168
rect 43 -175 52 -168
rect 32 -179 52 -175
rect 64 -179 68 -159
rect 18 -185 26 -179
rect 60 -185 68 -179
rect -18 -187 92 -185
rect -18 -199 -2 -187
rect 5 -199 23 -187
rect 30 -199 61 -187
rect 68 -199 92 -187
rect -18 -201 92 -199
<< metal2 >>
rect -5 241 1 279
rect 17 256 30 257
rect 17 250 23 256
rect 29 250 30 256
rect 17 249 30 250
rect 5 241 13 242
rect 11 235 13 241
rect 5 157 13 235
rect 17 169 25 249
rect 60 234 67 240
rect 35 213 36 219
rect 29 180 36 213
rect 29 175 44 180
rect 17 163 33 169
rect 5 151 9 157
rect 0 145 22 147
rect 0 138 15 145
rect 0 136 22 138
rect 0 -52 7 136
rect 27 111 33 163
rect 12 109 33 111
rect 18 103 33 109
rect 12 101 33 103
rect 37 97 44 175
rect 14 90 44 97
rect 14 58 23 90
rect 50 78 56 209
rect 60 159 66 234
rect 50 77 61 78
rect 51 71 54 77
rect 60 71 61 77
rect 51 70 61 71
rect 17 52 23 58
rect 14 -5 23 52
rect 70 34 76 209
rect 14 -11 16 -5
rect 22 -11 23 -5
rect 14 -13 23 -11
rect 37 32 76 34
rect 37 26 39 32
rect 45 26 76 32
rect 37 24 76 26
rect 37 -49 47 24
rect 23 -51 47 -49
rect 0 -54 19 -52
rect 0 -61 10 -54
rect 17 -61 19 -54
rect 23 -57 24 -51
rect 30 -57 47 -51
rect 23 -58 47 -57
rect 0 -63 19 -61
rect 46 -69 48 -63
rect 54 -69 56 -63
rect 2 -96 7 -90
rect -2 -148 7 -96
rect 4 -154 7 -148
rect 46 -147 56 -69
rect 46 -153 48 -147
rect 54 -153 56 -147
rect 46 -154 56 -153
rect 33 -168 46 -165
rect 33 -175 36 -168
rect 43 -175 46 -168
rect 33 -201 46 -175
<< ntransistor >>
rect 1 250 11 252
rect 54 250 64 252
rect 4 136 6 146
rect 56 136 58 146
rect 26 101 28 111
rect 64 101 66 111
rect 26 81 28 91
rect 64 81 66 91
rect 9 -73 19 -71
rect 9 -91 19 -89
rect 72 -79 74 -69
rect 72 -99 74 -89
rect 15 -141 17 -131
rect 57 -141 59 -131
<< ptransistor >>
rect 1 223 21 225
rect 44 223 64 225
rect 4 164 6 184
rect 56 164 58 184
rect 26 49 28 69
rect 64 49 66 69
rect 26 20 28 40
rect 64 20 66 40
rect 9 -24 29 -22
rect 9 -42 29 -40
rect 47 -43 49 -4
rect 72 -24 74 -4
rect 72 -53 74 -33
rect 15 -179 17 -159
rect 57 -179 59 -159
<< polycontact >>
rect 14 249 20 255
rect 32 221 38 227
rect 76 219 82 225
rect 41 209 47 215
rect -7 150 0 160
rect 36 150 43 160
rect 15 71 21 79
rect 28 72 40 78
rect 45 70 49 80
rect 74 73 79 79
rect 4 -11 12 -5
rect 58 -19 63 -8
rect 27 -71 32 -63
rect 58 -98 63 -90
rect 82 -98 88 -90
rect 25 -155 32 -145
rect 63 -155 70 -145
<< ndcontact >>
rect 1 253 11 257
rect 54 253 64 257
rect 1 245 11 249
rect 54 245 64 249
rect -1 136 3 146
rect 7 136 11 146
rect 51 136 55 146
rect 59 136 63 146
rect 21 101 25 111
rect 29 101 33 111
rect 59 101 63 111
rect 67 101 71 111
rect 21 81 25 91
rect 29 81 33 91
rect 59 81 63 91
rect 67 81 71 91
rect 9 -70 19 -66
rect 9 -78 19 -74
rect 9 -88 19 -84
rect 67 -79 71 -69
rect 75 -79 79 -69
rect 9 -96 19 -92
rect 67 -99 71 -89
rect 75 -99 79 -89
rect 10 -141 14 -131
rect 18 -141 22 -131
rect 52 -141 56 -131
rect 60 -141 64 -131
<< pdcontact >>
rect 1 226 21 230
rect 1 218 21 222
rect 44 226 64 230
rect 44 218 64 222
rect -1 164 3 184
rect 7 164 11 184
rect 51 164 55 184
rect 59 164 63 184
rect 21 49 25 69
rect 29 49 33 69
rect 59 49 63 69
rect 67 49 71 69
rect 21 20 25 40
rect 29 20 33 40
rect 59 20 63 40
rect 67 20 71 40
rect 9 -21 29 -17
rect 9 -29 29 -25
rect 9 -39 29 -35
rect 9 -47 29 -43
rect 42 -43 46 -4
rect 50 -43 54 -4
rect 67 -24 71 -4
rect 75 -24 79 -4
rect 67 -53 71 -33
rect 75 -53 79 -33
rect 10 -179 14 -159
rect 18 -179 22 -159
rect 52 -179 56 -159
rect 60 -179 64 -159
<< m2contact >>
rect 23 250 29 256
rect -5 235 1 241
rect 5 235 11 241
rect 67 234 73 240
rect 29 213 35 219
rect 50 209 56 215
rect 70 209 76 215
rect 9 151 15 157
rect 60 153 66 159
rect 15 138 22 145
rect 12 103 18 109
rect 11 52 17 58
rect 54 71 60 77
rect 39 26 45 32
rect 16 -11 22 -5
rect 10 -61 17 -54
rect 24 -57 30 -51
rect 48 -69 54 -63
rect -4 -96 2 -90
rect -2 -154 4 -148
rect 48 -153 54 -147
rect 36 -175 43 -168
<< psubstratepcontact >>
rect -4 265 3 277
rect 24 265 31 277
rect 53 265 60 277
rect -4 117 3 129
rect 24 117 31 129
rect 53 117 60 129
rect -4 -125 3 -113
rect 24 -125 31 -113
rect 53 -125 60 -113
<< nsubstratencontact >>
rect -2 191 5 203
rect 23 191 30 203
rect 61 191 68 203
rect -2 3 5 14
rect 23 3 30 14
rect 61 3 68 14
rect -2 -199 5 -187
rect 23 -199 30 -187
rect 61 -199 68 -187
<< labels >>
rlabel metal1 19 148 36 162 0 REGMEM
rlabel metal1 9 -84 42 -78 0 REGOUTn
rlabel polysilicon 46 42 51 70 0 INCLKLDn
rlabel metal1 36 32 59 40 0 INCLKn
rlabel metal1 79 73 92 79 0 CLKLD
rlabel polysilicon 82 91 92 99 0 CLK
rlabel metal1 -13 73 7 79 0 INCLKCLD
rlabel polysilicon -13 91 15 99 0 INCLK
rlabel metal2 33 -201 46 -175 0 REGOUT
rlabel polysilicon 82 -87 87 -67 0 RST
rlabel metal2 -5 241 1 279 0 REGIN
<< end >>
